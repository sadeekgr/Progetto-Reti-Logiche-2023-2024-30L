-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_12 is
end project_tb_12;

architecture project_tb_12_arch of project_tb_12 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    signal memory_control : std_logic := '0';

    -- first run
    constant SCENARIO_LENGTH : integer := 527;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;
    signal scenario_input : scenario_type := (121, 0, 171, 0, 244, 0, 11, 0, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 226, 0, 244, 0, 33, 0, 204, 0, 111, 0, 180, 0, 157, 0, 138, 0, 181, 0, 60, 0, 80, 0, 232, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 111, 0, 12, 0, 112, 0, 26, 0, 42, 0, 140, 0, 210, 0, 50, 0, 90, 0, 170, 0, 156, 0, 65, 0, 169, 0, 7, 0, 113, 0, 50, 0, 120, 0, 42, 0, 183, 0, 168, 0, 178, 0, 38, 0, 69, 0, 254, 0, 179, 0, 181, 0, 217, 0, 172, 0, 111, 0, 237, 0, 167, 0, 250, 0, 170, 0, 221, 0, 182, 0, 231, 0, 140, 0, 32, 0, 103, 0, 11, 0, 94, 0, 171, 0, 8, 0, 35, 0, 220, 0, 176, 0, 171, 0, 49, 0, 169, 0, 106, 0, 75, 0, 123, 0, 129, 0, 105, 0, 0, 0, 154, 0, 80, 0, 83, 0, 37, 0, 242, 0, 226, 0, 69, 0, 57, 0, 250, 0, 133, 0, 238, 0, 88, 0, 194, 0, 224, 0, 91, 0, 109, 0, 238, 0, 193, 0, 129, 0, 84, 0, 34, 0, 9, 0, 189, 0, 205, 0, 85, 0, 254, 0, 89, 0, 162, 0, 19, 0, 68, 0, 192, 0, 172, 0, 83, 0, 145, 0, 183, 0, 149, 0, 113, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 0, 71, 0, 19, 0, 14, 0, 178, 0, 53, 0, 126, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 249, 0, 253, 0, 140, 0, 208, 0, 127, 0, 139, 0, 221, 0, 219, 0, 31, 0, 13, 0, 148, 0, 128, 0, 105, 0, 45, 0, 20, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 249, 0, 136, 0, 68, 0, 10, 0, 226, 0, 11, 0, 121, 0, 245, 0, 150, 0, 136, 0, 69, 0, 64, 0, 224, 0, 136, 0, 197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 131, 0, 136, 0, 229, 0, 59, 0, 228, 0, 54, 0, 214, 0, 144, 0, 95, 0, 115, 0, 7, 0, 206, 0, 130, 0, 183, 0, 99, 0, 197, 0, 141, 0, 55, 0, 210, 0, 139, 0, 150, 0, 249, 0, 167, 0, 48, 0, 19, 0, 176, 0, 27, 0, 152, 0, 110, 0, 181, 0, 99, 0, 21, 0, 67, 0, 170, 0, 134, 0, 241, 0, 123, 0, 172, 0, 132, 0, 216, 0, 155, 0, 188, 0, 5, 0, 80, 0, 38, 0, 150, 0, 14, 0, 230, 0, 226, 0, 65, 0, 54, 0, 195, 0, 76, 0, 25, 0, 187, 0, 5, 0, 116, 0, 63, 0, 29, 0, 43, 0, 140, 0, 249, 0, 182, 0, 255, 0, 185, 0, 124, 0, 91, 0, 181, 0, 148, 0, 100, 0, 180, 0, 38, 0, 220, 0, 109, 0, 236, 0, 68, 0, 155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 99, 0, 236, 0, 71, 0, 230, 0, 159, 0, 30, 0, 159, 0, 239, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 179, 0, 114, 0, 192, 0, 14, 0, 58, 0, 221, 0, 9, 0, 172, 0, 152, 0, 103, 0, 32, 0, 245, 0, 210, 0, 241, 0, 243, 0, 128, 0, 172, 0, 39, 0, 69, 0, 224, 0, 232, 0, 179, 0, 72, 0, 177, 0, 84, 0, 216, 0, 148, 0, 183, 0, 240, 0, 202, 0, 98, 0, 32, 0, 248, 0, 42, 0, 56, 0, 165, 0, 252, 0, 14, 0, 97, 0, 174, 0, 80, 0, 103, 0, 213, 0, 141, 0, 163, 0, 67, 0, 188, 0, 6, 0, 100, 0, 101, 0, 205, 0, 19, 0, 159, 0, 148, 0);
    signal scenario_full  : scenario_type := (121, 31, 171, 31, 244, 31, 11, 31, 101, 31, 101, 30, 101, 29, 101, 28, 101, 27, 101, 26, 101, 25, 101, 24, 101, 23, 101, 22, 101, 21, 101, 20, 101, 19, 101, 18, 101, 17, 101, 16, 101, 15, 101, 14, 101, 13, 101, 12, 101, 11, 101, 10, 101, 9, 101, 8, 101, 7, 101, 6, 101, 5, 101, 4, 101, 3, 101, 2, 101, 1, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 101, 0, 226, 31, 244, 31, 33, 31, 204, 31, 111, 31, 180, 31, 157, 31, 138, 31, 181, 31, 60, 31, 80, 31, 232, 31, 232, 30, 232, 29, 232, 28, 232, 27, 232, 26, 232, 25, 232, 24, 232, 23, 232, 22, 232, 21, 232, 20, 232, 19, 232, 18, 232, 17, 232, 16, 40, 31, 111, 31, 12, 31, 112, 31, 26, 31, 42, 31, 140, 31, 210, 31, 50, 31, 90, 31, 170, 31, 156, 31, 65, 31, 169, 31, 7, 31, 113, 31, 50, 31, 120, 31, 42, 31, 183, 31, 168, 31, 178, 31, 38, 31, 69, 31, 254, 31, 179, 31, 181, 31, 217, 31, 172, 31, 111, 31, 237, 31, 167, 31, 250, 31, 170, 31, 221, 31, 182, 31, 231, 31, 140, 31, 32, 31, 103, 31, 11, 31, 94, 31, 171, 31, 8, 31, 35, 31, 220, 31, 176, 31, 171, 31, 49, 31, 169, 31, 106, 31, 75, 31, 123, 31, 129, 31, 105, 31, 105, 30, 154, 31, 80, 31, 83, 31, 37, 31, 242, 31, 226, 31, 69, 31, 57, 31, 250, 31, 133, 31, 238, 31, 88, 31, 194, 31, 224, 31, 91, 31, 109, 31, 238, 31, 193, 31, 129, 31, 84, 31, 34, 31, 9, 31, 189, 31, 205, 31, 85, 31, 254, 31, 89, 31, 162, 31, 19, 31, 68, 31, 192, 31, 172, 31, 83, 31, 145, 31, 183, 31, 149, 31, 113, 31, 113, 30, 113, 29, 113, 28, 113, 27, 113, 26, 113, 25, 113, 24, 113, 23, 113, 22, 113, 21, 113, 20, 113, 19, 113, 18, 113, 17, 78, 31, 71, 31, 19, 31, 14, 31, 178, 31, 53, 31, 126, 31, 126, 30, 126, 29, 126, 28, 126, 27, 126, 26, 126, 25, 126, 24, 126, 23, 126, 22, 126, 21, 126, 20, 126, 19, 126, 18, 126, 17, 249, 31, 253, 31, 140, 31, 208, 31, 127, 31, 139, 31, 221, 31, 219, 31, 31, 31, 13, 31, 148, 31, 128, 31, 105, 31, 45, 31, 20, 31, 41, 31, 41, 30, 41, 29, 41, 28, 41, 27, 41, 26, 41, 25, 41, 24, 41, 23, 41, 22, 41, 21, 41, 20, 41, 19, 41, 18, 41, 17, 41, 16, 41, 15, 41, 14, 41, 13, 249, 31, 136, 31, 68, 31, 10, 31, 226, 31, 11, 31, 121, 31, 245, 31, 150, 31, 136, 31, 69, 31, 64, 31, 224, 31, 136, 31, 197, 31, 197, 30, 197, 29, 197, 28, 197, 27, 197, 26, 197, 25, 197, 24, 197, 23, 197, 22, 197, 21, 197, 20, 197, 19, 197, 18, 197, 17, 197, 16, 197, 15, 197, 14, 197, 13, 197, 12, 197, 11, 197, 10, 197, 9, 197, 8, 197, 7, 197, 6, 197, 5, 197, 4, 6, 31, 131, 31, 136, 31, 229, 31, 59, 31, 228, 31, 54, 31, 214, 31, 144, 31, 95, 31, 115, 31, 7, 31, 206, 31, 130, 31, 183, 31, 99, 31, 197, 31, 141, 31, 55, 31, 210, 31, 139, 31, 150, 31, 249, 31, 167, 31, 48, 31, 19, 31, 176, 31, 27, 31, 152, 31, 110, 31, 181, 31, 99, 31, 21, 31, 67, 31, 170, 31, 134, 31, 241, 31, 123, 31, 172, 31, 132, 31, 216, 31, 155, 31, 188, 31, 5, 31, 80, 31, 38, 31, 150, 31, 14, 31, 230, 31, 226, 31, 65, 31, 54, 31, 195, 31, 76, 31, 25, 31, 187, 31, 5, 31, 116, 31, 63, 31, 29, 31, 43, 31, 140, 31, 249, 31, 182, 31, 255, 31, 185, 31, 124, 31, 91, 31, 181, 31, 148, 31, 100, 31, 180, 31, 38, 31, 220, 31, 109, 31, 236, 31, 68, 31, 155, 31, 155, 30, 155, 29, 155, 28, 155, 27, 155, 26, 155, 25, 155, 24, 155, 23, 155, 22, 155, 21, 155, 20, 155, 19, 155, 18, 155, 17, 155, 16, 155, 15, 155, 14, 155, 13, 155, 12, 155, 11, 155, 10, 155, 9, 155, 8, 155, 7, 155, 6, 155, 5, 155, 4, 155, 3, 155, 2, 155, 1, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 155, 0, 99, 31, 236, 31, 71, 31, 230, 31, 159, 31, 30, 31, 159, 31, 239, 31, 239, 30, 239, 29, 239, 28, 239, 27, 239, 26, 239, 25, 239, 24, 239, 23, 239, 22, 239, 21, 239, 20, 239, 19, 239, 18, 239, 17, 239, 16, 239, 15, 239, 14, 239, 13, 239, 12, 239, 11, 239, 10, 239, 9, 239, 8, 239, 7, 239, 6, 239, 5, 239, 4, 239, 3, 239, 2, 239, 1, 239, 0, 239, 0, 239, 0, 239, 0, 239, 0, 239, 0, 239, 0, 239, 0, 239, 0, 239, 0, 179, 31, 114, 31, 192, 31, 14, 31, 58, 31, 221, 31, 9, 31, 172, 31, 152, 31, 103, 31, 32, 31, 245, 31, 210, 31, 241, 31, 243, 31, 128, 31, 172, 31, 39, 31, 69, 31, 224, 31, 232, 31, 179, 31, 72, 31, 177, 31, 84, 31, 216, 31, 148, 31, 183, 31, 240, 31, 202, 31, 98, 31, 32, 31, 248, 31, 42, 31, 56, 31, 165, 31, 252, 31, 14, 31, 97, 31, 174, 31, 80, 31, 103, 31, 213, 31, 141, 31, 163, 31, 67, 31, 188, 31, 6, 31, 100, 31, 101, 31, 205, 31, 19, 31, 159, 31, 148, 31);
    constant SCENARIO_ADDRESS : integer := 890;

    -- second run

    constant SCENARIO_LENGTH_2 : integer := 252;
    type scenario_type_2 is array (0 to SCENARIO_LENGTH_2*2-1) of integer;
    signal scenario_input_2 : scenario_type_2 := (143, 0, 251, 0, 41, 0, 214, 0, 235, 0, 107, 0, 127, 0, 20, 0, 33, 0, 236, 0, 181, 0, 169, 0, 107, 0, 189, 0, 242, 0, 156, 0, 43, 0, 200, 0, 178, 0, 102, 0, 93, 0, 38, 0, 212, 0, 34, 0, 49, 0, 23, 0, 188, 0, 54, 0, 247, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 18, 0, 153, 0, 109, 0, 251, 0, 199, 0, 245, 0, 157, 0, 139, 0, 243, 0, 27, 0, 178, 0, 211, 0, 67, 0, 233, 0, 219, 0, 251, 0, 22, 0, 13, 0, 183, 0, 116, 0, 3, 0, 116, 0, 190, 0, 76, 0, 168, 0, 48, 0, 2, 0, 144, 0, 134, 0, 234, 0, 29, 0, 29, 0, 146, 0, 204, 0, 63, 0, 205, 0, 96, 0, 197, 0, 184, 0, 173, 0, 202, 0, 60, 0, 92, 0, 179, 0, 217, 0, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 189, 0, 75, 0, 55, 0, 202, 0, 48, 0, 93, 0, 0, 0, 0, 0, 0, 0, 200, 0, 155, 0, 126, 0, 42, 0, 107, 0, 164, 0, 254, 0, 36, 0, 180, 0, 87, 0, 182, 0, 150, 0, 135, 0, 188, 0, 200, 0, 78, 0, 164, 0, 124, 0, 55, 0, 249, 0, 241, 0, 93, 0, 99, 0, 8, 0, 180, 0, 56, 0, 215, 0, 145, 0, 88, 0, 138, 0, 107, 0, 74, 0, 93, 0, 244, 0, 4, 0, 120, 0, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 178, 0, 152, 0, 201, 0, 99, 0, 204, 0, 104, 0, 194, 0, 137, 0, 154, 0, 18, 0, 242, 0, 247, 0, 160, 0, 64, 0, 194, 0, 199, 0, 105, 0, 12, 0, 157, 0, 242, 0, 220, 0, 15, 0, 134, 0, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);
    signal scenario_full_2  : scenario_type_2 := (143, 31, 251, 31, 41, 31, 214, 31, 235, 31, 107, 31, 127, 31, 20, 31, 33, 31, 236, 31, 181, 31, 169, 31, 107, 31, 189, 31, 242, 31, 156, 31, 43, 31, 200, 31, 178, 31, 102, 31, 93, 31, 38, 31, 212, 31, 34, 31, 49, 31, 23, 31, 188, 31, 54, 31, 247, 31, 247, 30, 247, 29, 247, 28, 247, 27, 247, 26, 247, 25, 247, 24, 247, 23, 247, 22, 247, 21, 247, 20, 247, 19, 247, 18, 247, 17, 247, 16, 247, 15, 247, 14, 247, 13, 247, 12, 247, 11, 247, 10, 247, 9, 247, 8, 247, 7, 247, 6, 247, 5, 247, 4, 247, 3, 247, 2, 247, 1, 247, 0, 247, 0, 247, 0, 247, 0, 247, 0, 7, 31, 18, 31, 153, 31, 109, 31, 251, 31, 199, 31, 245, 31, 157, 31, 139, 31, 243, 31, 27, 31, 178, 31, 211, 31, 67, 31, 233, 31, 219, 31, 251, 31, 22, 31, 13, 31, 183, 31, 116, 31, 3, 31, 116, 31, 190, 31, 76, 31, 168, 31, 48, 31, 2, 31, 144, 31, 134, 31, 234, 31, 29, 31, 29, 31, 146, 31, 204, 31, 63, 31, 205, 31, 96, 31, 197, 31, 184, 31, 173, 31, 202, 31, 60, 31, 92, 31, 179, 31, 217, 31, 95, 31, 95, 30, 95, 29, 95, 28, 95, 27, 95, 26, 95, 25, 95, 24, 95, 23, 95, 22, 95, 21, 95, 20, 95, 19, 95, 18, 95, 17, 95, 16, 95, 15, 95, 14, 95, 13, 95, 12, 95, 11, 189, 31, 75, 31, 55, 31, 202, 31, 48, 31, 93, 31, 93, 30, 93, 29, 93, 28, 200, 31, 155, 31, 126, 31, 42, 31, 107, 31, 164, 31, 254, 31, 36, 31, 180, 31, 87, 31, 182, 31, 150, 31, 135, 31, 188, 31, 200, 31, 78, 31, 164, 31, 124, 31, 55, 31, 249, 31, 241, 31, 93, 31, 99, 31, 8, 31, 180, 31, 56, 31, 215, 31, 145, 31, 88, 31, 138, 31, 107, 31, 74, 31, 93, 31, 244, 31, 4, 31, 120, 31, 83, 31, 83, 30, 83, 29, 83, 28, 83, 27, 83, 26, 83, 25, 83, 24, 83, 23, 83, 22, 83, 21, 83, 20, 83, 19, 83, 18, 83, 17, 83, 16, 83, 15, 83, 14, 83, 13, 83, 12, 83, 11, 83, 10, 83, 9, 83, 8, 83, 7, 83, 6, 83, 5, 83, 4, 83, 3, 83, 2, 83, 1, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 83, 0, 20, 31, 178, 31, 152, 31, 201, 31, 99, 31, 204, 31, 104, 31, 194, 31, 137, 31, 154, 31, 18, 31, 242, 31, 247, 31, 160, 31, 64, 31, 194, 31, 199, 31, 105, 31, 12, 31, 157, 31, 242, 31, 220, 31, 15, 31, 134, 31, 102, 31, 102, 30, 102, 29, 102, 28, 102, 27, 102, 26, 102, 25);
    constant SCENARIO_ADDRESS_2 : integer := 10800;


    -- third run

    constant SCENARIO_LENGTH_3 : integer := 148;
    type scenario_type_3 is array (0 to SCENARIO_LENGTH_3*2-1) of integer;
    signal scenario_input_3 : scenario_type_3 := (160, 0, 95, 0, 92, 0, 134, 0, 226, 0, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 0, 98, 0, 157, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 231, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);
    signal scenario_full_3  : scenario_type_3 := (160, 31, 95, 31, 92, 31, 134, 31, 226, 31, 108, 31, 108, 30, 108, 29, 108, 28, 108, 27, 108, 26, 108, 25, 108, 24, 108, 23, 108, 22, 108, 21, 108, 20, 108, 19, 108, 18, 108, 17, 108, 16, 108, 15, 108, 14, 108, 13, 108, 12, 108, 11, 108, 10, 108, 9, 108, 8, 108, 7, 108, 6, 108, 5, 108, 4, 108, 3, 108, 2, 108, 1, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 108, 0, 80, 31, 98, 31, 157, 31, 157, 30, 157, 29, 157, 28, 157, 27, 157, 26, 157, 25, 157, 24, 157, 23, 157, 22, 157, 21, 157, 20, 157, 19, 157, 18, 157, 17, 157, 16, 157, 15, 157, 14, 157, 13, 157, 12, 157, 11, 157, 10, 157, 9, 157, 8, 157, 7, 157, 6, 157, 5, 157, 4, 157, 3, 157, 2, 157, 1, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 157, 0, 231, 31, 231, 30, 231, 29, 231, 28, 231, 27, 231, 26, 231, 25, 231, 24, 231, 23, 231, 22, 231, 21, 231, 20, 231, 19, 231, 18, 231, 17, 231, 16, 231, 15, 231, 14, 231, 13, 231, 12, 231, 11, 231, 10, 231, 9, 231, 8, 231, 7, 231, 6, 231, 5, 231, 4, 231, 3, 231, 2, 231, 1, 231, 0, 231, 0, 231, 0, 231, 0);
    constant SCENARIO_ADDRESS_3 : integer := 21610;


    -- fourth run
    
    constant SCENARIO_LENGTH_4 : integer := 709;
    type scenario_type_4 is array (0 to SCENARIO_LENGTH_4*2-1) of integer;
    signal scenario_input_4 : scenario_type_4 := (248, 0, 18, 0, 45, 0, 90, 0, 119, 0, 224, 0, 102, 0, 227, 0, 129, 0, 76, 0, 141, 0, 220, 0, 21, 0, 55, 0, 156, 0, 126, 0, 75, 0, 34, 0, 155, 0, 91, 0, 28, 0, 162, 0, 95, 0, 207, 0, 184, 0, 19, 0, 66, 0, 101, 0, 49, 0, 188, 0, 78, 0, 167, 0, 163, 0, 57, 0, 41, 0, 60, 0, 194, 0, 211, 0, 14, 0, 157, 0, 30, 0, 201, 0, 245, 0, 180, 0, 112, 0, 121, 0, 213, 0, 179, 0, 41, 0, 76, 0, 176, 0, 209, 0, 161, 0, 139, 0, 203, 0, 211, 0, 216, 0, 106, 0, 112, 0, 19, 0, 119, 0, 26, 0, 121, 0, 97, 0, 15, 0, 45, 0, 212, 0, 222, 0, 244, 0, 189, 0, 6, 0, 96, 0, 70, 0, 5, 0, 34, 0, 212, 0, 189, 0, 209, 0, 148, 0, 53, 0, 130, 0, 219, 0, 145, 0, 141, 0, 190, 0, 79, 0, 6, 0, 201, 0, 162, 0, 84, 0, 90, 0, 121, 0, 167, 0, 186, 0, 229, 0, 155, 0, 21, 0, 167, 0, 160, 0, 149, 0, 182, 0, 144, 0, 135, 0, 140, 0, 209, 0, 236, 0, 7, 0, 177, 0, 131, 0, 135, 0, 107, 0, 225, 0, 214, 0, 100, 0, 195, 0, 138, 0, 154, 0, 94, 0, 226, 0, 8, 0, 7, 0, 179, 0, 184, 0, 89, 0, 123, 0, 139, 0, 220, 0, 20, 0, 105, 0, 169, 0, 139, 0, 132, 0, 21, 0, 205, 0, 136, 0, 112, 0, 100, 0, 182, 0, 45, 0, 222, 0, 228, 0, 171, 0, 30, 0, 104, 0, 115, 0, 14, 0, 231, 0, 111, 0, 161, 0, 102, 0, 213, 0, 76, 0, 28, 0, 134, 0, 99, 0, 122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 233, 0, 231, 0, 255, 0, 243, 0, 130, 0, 106, 0, 196, 0, 110, 0, 88, 0, 138, 0, 165, 0, 110, 0, 19, 0, 12, 0, 228, 0, 210, 0, 152, 0, 170, 0, 163, 0, 199, 0, 74, 0, 230, 0, 46, 0, 231, 0, 116, 0, 173, 0, 185, 0, 32, 0, 249, 0, 132, 0, 213, 0, 73, 0, 210, 0, 235, 0, 13, 0, 29, 0, 165, 0, 254, 0, 189, 0, 139, 0, 155, 0, 50, 0, 14, 0, 153, 0, 72, 0, 20, 0, 50, 0, 195, 0, 236, 0, 243, 0, 238, 0, 217, 0, 126, 0, 95, 0, 184, 0, 219, 0, 76, 0, 19, 0, 44, 0, 195, 0, 230, 0, 0, 0, 38, 0, 85, 0, 59, 0, 90, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 99, 0, 50, 0, 81, 0, 91, 0, 51, 0, 161, 0, 115, 0, 81, 0, 75, 0, 228, 0, 107, 0, 145, 0, 109, 0, 186, 0, 145, 0, 209, 0, 49, 0, 244, 0, 38, 0, 178, 0, 48, 0, 148, 0, 15, 0, 250, 0, 115, 0, 153, 0, 84, 0, 173, 0, 206, 0, 242, 0, 145, 0, 120, 0, 255, 0, 227, 0, 82, 0, 245, 0, 103, 0, 227, 0, 195, 0, 249, 0, 77, 0, 86, 0, 123, 0, 247, 0, 42, 0, 40, 0, 6, 0, 2, 0, 213, 0, 70, 0, 18, 0, 140, 0, 19, 0, 132, 0, 6, 0, 119, 0, 211, 0, 168, 0, 210, 0, 196, 0, 97, 0, 224, 0, 49, 0, 14, 0, 24, 0, 220, 0, 110, 0, 204, 0, 255, 0, 39, 0, 20, 0, 231, 0, 153, 0, 50, 0, 246, 0, 125, 0, 173, 0, 153, 0, 51, 0, 238, 0, 209, 0, 120, 0, 53, 0, 253, 0, 188, 0, 213, 0, 123, 0, 183, 0, 113, 0, 19, 0, 54, 0, 215, 0, 139, 0, 51, 0, 134, 0, 220, 0, 173, 0, 40, 0, 152, 0, 133, 0, 224, 0, 76, 0, 254, 0, 39, 0, 147, 0, 225, 0, 108, 0, 160, 0, 114, 0, 214, 0, 57, 0, 24, 0, 13, 0, 136, 0, 207, 0, 3, 0, 132, 0, 25, 0, 111, 0, 136, 0, 131, 0, 191, 0, 27, 0, 25, 0, 189, 0, 100, 0, 180, 0, 70, 0, 72, 0, 227, 0, 172, 0, 33, 0, 59, 0, 27, 0, 112, 0, 116, 0, 178, 0, 128, 0, 105, 0, 216, 0, 250, 0, 231, 0, 92, 0, 218, 0, 124, 0, 179, 0, 9, 0, 94, 0, 140, 0, 15, 0, 212, 0, 213, 0, 15, 0, 2, 0, 124, 0, 223, 0, 66, 0, 226, 0, 173, 0, 92, 0, 245, 0, 77, 0, 4, 0, 12, 0, 208, 0, 6, 0, 183, 0, 221, 0, 234, 0, 240, 0, 139, 0, 176, 0, 15, 0, 172, 0, 80, 0, 224, 0, 88, 0, 212, 0, 27, 0, 15, 0, 54, 0, 166, 0, 84, 0, 128, 0, 250, 0, 254, 0, 24, 0, 158, 0, 121, 0, 13, 0, 246, 0, 35, 0, 116, 0, 235, 0, 13, 0, 191, 0, 136, 0, 143, 0, 150, 0, 225, 0, 136, 0, 250, 0, 152, 0, 187, 0, 31, 0, 89, 0, 63, 0, 15, 0, 110, 0, 53, 0, 21, 0, 254, 0, 68, 0, 197, 0, 115, 0, 238, 0, 32, 0, 213, 0, 128, 0, 164, 0, 201, 0, 38, 0, 182, 0, 73, 0, 35, 0, 12, 0, 169, 0, 104, 0, 116, 0, 210, 0, 181, 0, 207, 0, 227, 0, 215, 0, 153, 0, 118, 0, 25, 0, 17, 0, 56, 0, 66, 0, 234, 0, 247, 0, 238, 0, 68, 0, 120, 0, 136, 0, 194, 0, 188, 0, 95, 0, 141, 0, 181, 0, 144, 0, 165, 0, 187, 0, 161, 0, 40, 0, 131, 0, 252, 0, 179, 0, 210, 0, 239, 0, 223, 0, 251, 0, 169, 0, 51, 0, 142, 0, 91, 0, 64, 0, 6, 0, 28, 0, 201, 0, 34, 0, 12, 0, 177, 0, 224, 0, 219, 0, 22, 0, 170, 0, 43, 0, 56, 0, 182, 0, 158, 0, 250, 0, 186, 0, 181, 0, 44, 0, 197, 0, 178, 0, 73, 0, 224, 0, 140, 0, 173, 0, 54, 0, 231, 0, 152, 0, 22, 0, 253, 0, 196, 0, 219, 0, 12, 0, 188, 0, 219, 0, 31, 0, 137, 0, 8, 0, 17, 0, 222, 0, 182, 0, 163, 0, 248, 0, 226, 0, 98, 0, 231, 0, 191, 0, 2, 0, 9, 0, 244, 0, 200, 0, 140, 0, 107, 0, 97, 0, 7, 0, 31, 0, 37, 0, 40, 0, 87, 0, 26, 0, 148, 0, 41, 0, 27, 0, 208, 0, 174, 0, 120, 0, 68, 0, 21, 0, 15, 0, 200, 0, 127, 0, 93, 0, 12, 0, 80, 0, 131, 0, 247, 0, 7, 0, 215, 0, 189, 0, 215, 0, 188, 0, 213, 0, 84, 0, 112, 0, 77, 0, 144, 0, 81, 0, 101, 0, 196, 0, 26, 0, 82, 0, 174, 0, 170, 0, 186, 0, 49, 0, 244, 0, 115, 0, 218, 0, 6, 0, 49, 0, 20, 0, 46, 0, 126, 0, 186, 0, 84, 0, 67, 0, 11, 0, 105, 0, 100, 0, 102, 0, 136, 0, 237, 0, 200, 0, 203, 0, 177, 0, 55, 0, 204, 0, 209, 0, 208, 0, 108, 0, 15, 0, 30, 0, 240, 0, 13, 0, 191, 0, 125, 0, 88, 0, 193, 0, 192, 0, 124, 0, 53, 0, 82, 0, 93, 0, 95, 0, 90, 0, 25, 0, 132, 0, 209, 0, 155, 0, 125, 0, 236, 0, 92, 0, 236, 0, 29, 0, 61, 0, 94, 0, 42, 0, 133, 0, 52, 0, 114, 0, 173, 0, 182, 0, 240, 0, 33, 0, 102, 0, 207, 0, 28, 0, 26, 0, 27, 0, 59, 0, 250, 0, 59, 0, 70, 0, 148, 0, 143, 0, 242, 0, 96, 0, 149, 0, 45, 0, 111, 0, 151, 0, 248, 0, 145, 0, 106, 0, 168, 0, 107, 0, 9, 0, 18, 0, 178, 0, 196, 0, 179, 0, 141, 0, 165, 0, 185, 0, 4, 0, 204, 0, 122, 0, 6, 0, 230, 0, 105, 0, 22, 0, 102, 0, 172, 0, 248, 0, 196, 0, 70, 0, 184, 0, 114, 0, 169, 0, 239, 0, 9, 0, 0, 0, 0, 0, 0, 0);
    signal scenario_full_4  : scenario_type_4 := (248, 31, 18, 31, 45, 31, 90, 31, 119, 31, 224, 31, 102, 31, 227, 31, 129, 31, 76, 31, 141, 31, 220, 31, 21, 31, 55, 31, 156, 31, 126, 31, 75, 31, 34, 31, 155, 31, 91, 31, 28, 31, 162, 31, 95, 31, 207, 31, 184, 31, 19, 31, 66, 31, 101, 31, 49, 31, 188, 31, 78, 31, 167, 31, 163, 31, 57, 31, 41, 31, 60, 31, 194, 31, 211, 31, 14, 31, 157, 31, 30, 31, 201, 31, 245, 31, 180, 31, 112, 31, 121, 31, 213, 31, 179, 31, 41, 31, 76, 31, 176, 31, 209, 31, 161, 31, 139, 31, 203, 31, 211, 31, 216, 31, 106, 31, 112, 31, 19, 31, 119, 31, 26, 31, 121, 31, 97, 31, 15, 31, 45, 31, 212, 31, 222, 31, 244, 31, 189, 31, 6, 31, 96, 31, 70, 31, 5, 31, 34, 31, 212, 31, 189, 31, 209, 31, 148, 31, 53, 31, 130, 31, 219, 31, 145, 31, 141, 31, 190, 31, 79, 31, 6, 31, 201, 31, 162, 31, 84, 31, 90, 31, 121, 31, 167, 31, 186, 31, 229, 31, 155, 31, 21, 31, 167, 31, 160, 31, 149, 31, 182, 31, 144, 31, 135, 31, 140, 31, 209, 31, 236, 31, 7, 31, 177, 31, 131, 31, 135, 31, 107, 31, 225, 31, 214, 31, 100, 31, 195, 31, 138, 31, 154, 31, 94, 31, 226, 31, 8, 31, 7, 31, 179, 31, 184, 31, 89, 31, 123, 31, 139, 31, 220, 31, 20, 31, 105, 31, 169, 31, 139, 31, 132, 31, 21, 31, 205, 31, 136, 31, 112, 31, 100, 31, 182, 31, 45, 31, 222, 31, 228, 31, 171, 31, 30, 31, 104, 31, 115, 31, 14, 31, 231, 31, 111, 31, 161, 31, 102, 31, 213, 31, 76, 31, 28, 31, 134, 31, 99, 31, 122, 31, 122, 30, 122, 29, 122, 28, 122, 27, 122, 26, 122, 25, 122, 24, 122, 23, 122, 22, 122, 21, 122, 20, 233, 31, 231, 31, 255, 31, 243, 31, 130, 31, 106, 31, 196, 31, 110, 31, 88, 31, 138, 31, 165, 31, 110, 31, 19, 31, 12, 31, 228, 31, 210, 31, 152, 31, 170, 31, 163, 31, 199, 31, 74, 31, 230, 31, 46, 31, 231, 31, 116, 31, 173, 31, 185, 31, 32, 31, 249, 31, 132, 31, 213, 31, 73, 31, 210, 31, 235, 31, 13, 31, 29, 31, 165, 31, 254, 31, 189, 31, 139, 31, 155, 31, 50, 31, 14, 31, 153, 31, 72, 31, 20, 31, 50, 31, 195, 31, 236, 31, 243, 31, 238, 31, 217, 31, 126, 31, 95, 31, 184, 31, 219, 31, 76, 31, 19, 31, 44, 31, 195, 31, 230, 31, 230, 30, 38, 31, 85, 31, 59, 31, 90, 31, 84, 31, 84, 30, 84, 29, 84, 28, 84, 27, 99, 31, 50, 31, 81, 31, 91, 31, 51, 31, 161, 31, 115, 31, 81, 31, 75, 31, 228, 31, 107, 31, 145, 31, 109, 31, 186, 31, 145, 31, 209, 31, 49, 31, 244, 31, 38, 31, 178, 31, 48, 31, 148, 31, 15, 31, 250, 31, 115, 31, 153, 31, 84, 31, 173, 31, 206, 31, 242, 31, 145, 31, 120, 31, 255, 31, 227, 31, 82, 31, 245, 31, 103, 31, 227, 31, 195, 31, 249, 31, 77, 31, 86, 31, 123, 31, 247, 31, 42, 31, 40, 31, 6, 31, 2, 31, 213, 31, 70, 31, 18, 31, 140, 31, 19, 31, 132, 31, 6, 31, 119, 31, 211, 31, 168, 31, 210, 31, 196, 31, 97, 31, 224, 31, 49, 31, 14, 31, 24, 31, 220, 31, 110, 31, 204, 31, 255, 31, 39, 31, 20, 31, 231, 31, 153, 31, 50, 31, 246, 31, 125, 31, 173, 31, 153, 31, 51, 31, 238, 31, 209, 31, 120, 31, 53, 31, 253, 31, 188, 31, 213, 31, 123, 31, 183, 31, 113, 31, 19, 31, 54, 31, 215, 31, 139, 31, 51, 31, 134, 31, 220, 31, 173, 31, 40, 31, 152, 31, 133, 31, 224, 31, 76, 31, 254, 31, 39, 31, 147, 31, 225, 31, 108, 31, 160, 31, 114, 31, 214, 31, 57, 31, 24, 31, 13, 31, 136, 31, 207, 31, 3, 31, 132, 31, 25, 31, 111, 31, 136, 31, 131, 31, 191, 31, 27, 31, 25, 31, 189, 31, 100, 31, 180, 31, 70, 31, 72, 31, 227, 31, 172, 31, 33, 31, 59, 31, 27, 31, 112, 31, 116, 31, 178, 31, 128, 31, 105, 31, 216, 31, 250, 31, 231, 31, 92, 31, 218, 31, 124, 31, 179, 31, 9, 31, 94, 31, 140, 31, 15, 31, 212, 31, 213, 31, 15, 31, 2, 31, 124, 31, 223, 31, 66, 31, 226, 31, 173, 31, 92, 31, 245, 31, 77, 31, 4, 31, 12, 31, 208, 31, 6, 31, 183, 31, 221, 31, 234, 31, 240, 31, 139, 31, 176, 31, 15, 31, 172, 31, 80, 31, 224, 31, 88, 31, 212, 31, 27, 31, 15, 31, 54, 31, 166, 31, 84, 31, 128, 31, 250, 31, 254, 31, 24, 31, 158, 31, 121, 31, 13, 31, 246, 31, 35, 31, 116, 31, 235, 31, 13, 31, 191, 31, 136, 31, 143, 31, 150, 31, 225, 31, 136, 31, 250, 31, 152, 31, 187, 31, 31, 31, 89, 31, 63, 31, 15, 31, 110, 31, 53, 31, 21, 31, 254, 31, 68, 31, 197, 31, 115, 31, 238, 31, 32, 31, 213, 31, 128, 31, 164, 31, 201, 31, 38, 31, 182, 31, 73, 31, 35, 31, 12, 31, 169, 31, 104, 31, 116, 31, 210, 31, 181, 31, 207, 31, 227, 31, 215, 31, 153, 31, 118, 31, 25, 31, 17, 31, 56, 31, 66, 31, 234, 31, 247, 31, 238, 31, 68, 31, 120, 31, 136, 31, 194, 31, 188, 31, 95, 31, 141, 31, 181, 31, 144, 31, 165, 31, 187, 31, 161, 31, 40, 31, 131, 31, 252, 31, 179, 31, 210, 31, 239, 31, 223, 31, 251, 31, 169, 31, 51, 31, 142, 31, 91, 31, 64, 31, 6, 31, 28, 31, 201, 31, 34, 31, 12, 31, 177, 31, 224, 31, 219, 31, 22, 31, 170, 31, 43, 31, 56, 31, 182, 31, 158, 31, 250, 31, 186, 31, 181, 31, 44, 31, 197, 31, 178, 31, 73, 31, 224, 31, 140, 31, 173, 31, 54, 31, 231, 31, 152, 31, 22, 31, 253, 31, 196, 31, 219, 31, 12, 31, 188, 31, 219, 31, 31, 31, 137, 31, 8, 31, 17, 31, 222, 31, 182, 31, 163, 31, 248, 31, 226, 31, 98, 31, 231, 31, 191, 31, 2, 31, 9, 31, 244, 31, 200, 31, 140, 31, 107, 31, 97, 31, 7, 31, 31, 31, 37, 31, 40, 31, 87, 31, 26, 31, 148, 31, 41, 31, 27, 31, 208, 31, 174, 31, 120, 31, 68, 31, 21, 31, 15, 31, 200, 31, 127, 31, 93, 31, 12, 31, 80, 31, 131, 31, 247, 31, 7, 31, 215, 31, 189, 31, 215, 31, 188, 31, 213, 31, 84, 31, 112, 31, 77, 31, 144, 31, 81, 31, 101, 31, 196, 31, 26, 31, 82, 31, 174, 31, 170, 31, 186, 31, 49, 31, 244, 31, 115, 31, 218, 31, 6, 31, 49, 31, 20, 31, 46, 31, 126, 31, 186, 31, 84, 31, 67, 31, 11, 31, 105, 31, 100, 31, 102, 31, 136, 31, 237, 31, 200, 31, 203, 31, 177, 31, 55, 31, 204, 31, 209, 31, 208, 31, 108, 31, 15, 31, 30, 31, 240, 31, 13, 31, 191, 31, 125, 31, 88, 31, 193, 31, 192, 31, 124, 31, 53, 31, 82, 31, 93, 31, 95, 31, 90, 31, 25, 31, 132, 31, 209, 31, 155, 31, 125, 31, 236, 31, 92, 31, 236, 31, 29, 31, 61, 31, 94, 31, 42, 31, 133, 31, 52, 31, 114, 31, 173, 31, 182, 31, 240, 31, 33, 31, 102, 31, 207, 31, 28, 31, 26, 31, 27, 31, 59, 31, 250, 31, 59, 31, 70, 31, 148, 31, 143, 31, 242, 31, 96, 31, 149, 31, 45, 31, 111, 31, 151, 31, 248, 31, 145, 31, 106, 31, 168, 31, 107, 31, 9, 31, 18, 31, 178, 31, 196, 31, 179, 31, 141, 31, 165, 31, 185, 31, 4, 31, 204, 31, 122, 31, 6, 31, 230, 31, 105, 31, 22, 31, 102, 31, 172, 31, 248, 31, 196, 31, 70, 31, 184, 31, 114, 31, 169, 31, 239, 31, 9, 31, 9, 30, 9, 29, 9, 28);
    constant SCENARIO_ADDRESS_4 : integer := 31005;


    -- fifth run

    constant SCENARIO_LENGTH_5 : integer := 917;
    type scenario_type_5 is array (0 to SCENARIO_LENGTH_5*2-1) of integer;
    signal scenario_input_5 : scenario_type_5 := (54, 0, 180, 0, 150, 0, 177, 0, 76, 0, 67, 0, 152, 0, 218, 0, 190, 0, 184, 0, 172, 0, 3, 0, 148, 0, 189, 0, 251, 0, 220, 0, 164, 0, 3, 0, 194, 0, 204, 0, 141, 0, 108, 0, 127, 0, 87, 0, 199, 0, 160, 0, 20, 0, 19, 0, 242, 0, 133, 0, 195, 0, 12, 0, 78, 0, 59, 0, 56, 0, 227, 0, 20, 0, 145, 0, 237, 0, 131, 0, 11, 0, 121, 0, 117, 0, 239, 0, 157, 0, 111, 0, 131, 0, 10, 0, 172, 0, 234, 0, 196, 0, 101, 0, 146, 0, 177, 0, 1, 0, 38, 0, 51, 0, 80, 0, 199, 0, 89, 0, 91, 0, 123, 0, 20, 0, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 0, 241, 0, 92, 0, 140, 0, 221, 0, 243, 0, 94, 0, 21, 0, 46, 0, 50, 0, 192, 0, 147, 0, 5, 0, 153, 0, 243, 0, 150, 0, 229, 0, 231, 0, 31, 0, 229, 0, 31, 0, 24, 0, 254, 0, 215, 0, 124, 0, 40, 0, 137, 0, 0, 0, 56, 0, 199, 0, 253, 0, 52, 0, 17, 0, 206, 0, 146, 0, 219, 0, 206, 0, 5, 0, 56, 0, 58, 0, 175, 0, 104, 0, 186, 0, 172, 0, 202, 0, 177, 0, 28, 0, 208, 0, 145, 0, 214, 0, 1, 0, 177, 0, 7, 0, 28, 0, 103, 0, 155, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 237, 0, 99, 0, 133, 0, 184, 0, 215, 0, 240, 0, 247, 0, 109, 0, 200, 0, 97, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 150, 0, 148, 0, 220, 0, 31, 0, 103, 0, 144, 0, 178, 0, 236, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 162, 0, 121, 0, 199, 0, 149, 0, 167, 0, 45, 0, 254, 0, 154, 0, 163, 0, 146, 0, 34, 0, 190, 0, 155, 0, 241, 0, 143, 0, 34, 0, 165, 0, 58, 0, 17, 0, 44, 0, 63, 0, 70, 0, 164, 0, 47, 0, 3, 0, 236, 0, 177, 0, 158, 0, 220, 0, 179, 0, 1, 0, 240, 0, 218, 0, 139, 0, 149, 0, 166, 0, 243, 0, 208, 0, 123, 0, 140, 0, 8, 0, 66, 0, 51, 0, 162, 0, 135, 0, 19, 0, 143, 0, 172, 0, 248, 0, 16, 0, 77, 0, 103, 0, 102, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 219, 0, 196, 0, 25, 0, 2, 0, 163, 0, 204, 0, 125, 0, 50, 0, 56, 0, 206, 0, 70, 0, 32, 0, 32, 0, 61, 0, 158, 0, 56, 0, 166, 0, 223, 0, 111, 0, 95, 0, 83, 0, 225, 0, 229, 0, 84, 0, 134, 0, 94, 0, 9, 0, 53, 0, 129, 0, 119, 0, 118, 0, 244, 0, 250, 0, 159, 0, 190, 0, 200, 0, 115, 0, 134, 0, 72, 0, 205, 0, 105, 0, 154, 0, 168, 0, 133, 0, 109, 0, 185, 0, 54, 0, 36, 0, 121, 0, 26, 0, 74, 0, 4, 0, 13, 0, 250, 0, 77, 0, 151, 0, 28, 0, 113, 0, 194, 0, 56, 0, 81, 0, 51, 0, 131, 0, 21, 0, 162, 0, 121, 0, 125, 0, 212, 0, 255, 0, 123, 0, 163, 0, 102, 0, 253, 0, 76, 0, 201, 0, 233, 0, 232, 0, 178, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78, 0, 87, 0, 44, 0, 220, 0, 157, 0, 81, 0, 180, 0, 174, 0, 38, 0, 89, 0, 234, 0, 109, 0, 122, 0, 3, 0, 41, 0, 214, 0, 162, 0, 123, 0, 94, 0, 220, 0, 107, 0, 1, 0, 26, 0, 187, 0, 97, 0, 13, 0, 238, 0, 163, 0, 6, 0, 119, 0, 31, 0, 20, 0, 161, 0, 218, 0, 130, 0, 43, 0, 254, 0, 145, 0, 247, 0, 6, 0, 200, 0, 30, 0, 13, 0, 81, 0, 101, 0, 205, 0, 12, 0, 201, 0, 255, 0, 11, 0, 234, 0, 90, 0, 201, 0, 253, 0, 211, 0, 72, 0, 23, 0, 98, 0, 23, 0, 182, 0, 243, 0, 74, 0, 239, 0, 239, 0, 147, 0, 180, 0, 140, 0, 239, 0, 66, 0, 181, 0, 42, 0, 219, 0, 24, 0, 70, 0, 234, 0, 92, 0, 145, 0, 143, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 212, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 105, 0, 251, 0, 85, 0, 88, 0, 23, 0, 50, 0, 112, 0, 63, 0, 42, 0, 116, 0, 142, 0, 214, 0, 66, 0, 52, 0, 141, 0, 191, 0, 82, 0, 40, 0, 178, 0, 161, 0, 91, 0, 218, 0, 159, 0, 92, 0, 93, 0, 179, 0, 111, 0, 102, 0, 116, 0, 29, 0, 63, 0, 96, 0, 200, 0, 49, 0, 58, 0, 182, 0, 37, 0, 93, 0, 134, 0, 6, 0, 172, 0, 124, 0, 191, 0, 117, 0, 143, 0, 172, 0, 249, 0, 30, 0, 69, 0, 203, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 133, 0, 202, 0, 92, 0, 23, 0, 23, 0, 226, 0, 26, 0, 215, 0, 12, 0, 235, 0, 102, 0, 205, 0, 146, 0, 141, 0, 48, 0, 156, 0, 169, 0, 16, 0, 130, 0, 138, 0, 62, 0, 146, 0, 185, 0, 1, 0, 181, 0, 8, 0, 121, 0, 156, 0, 5, 0, 80, 0, 167, 0, 255, 0, 134, 0, 57, 0, 66, 0, 247, 0, 48, 0, 213, 0, 9, 0, 55, 0, 55, 0, 6, 0, 235, 0, 230, 0, 18, 0, 31, 0, 62, 0, 145, 0, 107, 0, 129, 0, 167, 0, 206, 0, 143, 0, 222, 0, 125, 0, 123, 0, 157, 0, 155, 0, 199, 0, 49, 0, 141, 0, 255, 0, 26, 0, 35, 0, 37, 0, 244, 0, 35, 0, 115, 0, 122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 208, 0, 74, 0, 116, 0, 177, 0, 228, 0, 44, 0, 200, 0, 255, 0, 134, 0, 108, 0, 35, 0, 194, 0, 223, 0, 119, 0, 105, 0, 30, 0, 35, 0, 196, 0, 157, 0, 109, 0, 209, 0, 204, 0, 0, 0, 79, 0, 17, 0, 201, 0, 253, 0, 46, 0, 131, 0, 131, 0, 252, 0, 122, 0, 200, 0, 159, 0, 193, 0, 10, 0, 196, 0, 139, 0, 224, 0, 210, 0, 2, 0, 212, 0, 153, 0, 32, 0, 225, 0, 33, 0, 8, 0, 5, 0, 245, 0, 152, 0, 132, 0, 28, 0, 66, 0, 60, 0, 213, 0, 127, 0, 14, 0, 101, 0, 172, 0, 124, 0, 91, 0, 154, 0, 194, 0, 193, 0, 22, 0, 127, 0, 110, 0, 49, 0, 179, 0, 22, 0, 135, 0, 119, 0, 141, 0, 97, 0, 64, 0, 23, 0, 56, 0, 144, 0, 221, 0, 12, 0, 244, 0, 61, 0, 65, 0, 156, 0, 102, 0, 228, 0, 195, 0, 35, 0, 32, 0, 206, 0, 57, 0, 129, 0, 148, 0, 38, 0, 89, 0, 89, 0, 239, 0, 191, 0, 165, 0, 73, 0, 64, 0, 128, 0, 155, 0, 41, 0, 217, 0, 195, 0, 221, 0, 31, 0, 181, 0, 160, 0, 161, 0, 41, 0, 144, 0, 128, 0, 236, 0, 46, 0, 163, 0, 69, 0, 50, 0, 9, 0, 171, 0, 239, 0, 186, 0, 57, 0, 192, 0, 197, 0, 176, 0, 2, 0, 157, 0, 200, 0, 90, 0, 76, 0, 52, 0);
    signal scenario_full_5  : scenario_type_5 := (54, 31, 180, 31, 150, 31, 177, 31, 76, 31, 67, 31, 152, 31, 218, 31, 190, 31, 184, 31, 172, 31, 3, 31, 148, 31, 189, 31, 251, 31, 220, 31, 164, 31, 3, 31, 194, 31, 204, 31, 141, 31, 108, 31, 127, 31, 87, 31, 199, 31, 160, 31, 20, 31, 19, 31, 242, 31, 133, 31, 195, 31, 12, 31, 78, 31, 59, 31, 56, 31, 227, 31, 20, 31, 145, 31, 237, 31, 131, 31, 11, 31, 121, 31, 117, 31, 239, 31, 157, 31, 111, 31, 131, 31, 10, 31, 172, 31, 234, 31, 196, 31, 101, 31, 146, 31, 177, 31, 1, 31, 38, 31, 51, 31, 80, 31, 199, 31, 89, 31, 91, 31, 123, 31, 20, 31, 73, 31, 73, 30, 73, 29, 73, 28, 73, 27, 73, 26, 73, 25, 73, 24, 73, 23, 73, 22, 73, 21, 73, 20, 73, 19, 73, 18, 73, 17, 73, 16, 73, 15, 73, 14, 73, 13, 73, 12, 73, 11, 73, 10, 73, 9, 73, 8, 73, 7, 73, 6, 73, 5, 73, 4, 60, 31, 241, 31, 92, 31, 140, 31, 221, 31, 243, 31, 94, 31, 21, 31, 46, 31, 50, 31, 192, 31, 147, 31, 5, 31, 153, 31, 243, 31, 150, 31, 229, 31, 231, 31, 31, 31, 229, 31, 31, 31, 24, 31, 254, 31, 215, 31, 124, 31, 40, 31, 137, 31, 137, 30, 56, 31, 199, 31, 253, 31, 52, 31, 17, 31, 206, 31, 146, 31, 219, 31, 206, 31, 5, 31, 56, 31, 58, 31, 175, 31, 104, 31, 186, 31, 172, 31, 202, 31, 177, 31, 28, 31, 208, 31, 145, 31, 214, 31, 1, 31, 177, 31, 7, 31, 28, 31, 103, 31, 155, 31, 155, 30, 155, 29, 155, 28, 155, 27, 155, 26, 155, 25, 155, 24, 155, 23, 155, 22, 155, 21, 155, 20, 155, 19, 155, 18, 155, 17, 155, 16, 155, 15, 155, 14, 155, 13, 155, 12, 155, 11, 155, 10, 155, 9, 155, 8, 155, 7, 155, 6, 155, 5, 155, 4, 155, 3, 170, 31, 237, 31, 99, 31, 133, 31, 184, 31, 215, 31, 240, 31, 247, 31, 109, 31, 200, 31, 97, 31, 97, 30, 97, 29, 97, 28, 97, 27, 97, 26, 97, 25, 97, 24, 97, 23, 97, 22, 97, 21, 97, 20, 97, 19, 97, 18, 97, 17, 97, 16, 97, 15, 97, 14, 97, 13, 97, 12, 97, 11, 97, 10, 97, 9, 97, 8, 97, 7, 97, 6, 97, 5, 97, 4, 97, 3, 97, 2, 33, 31, 150, 31, 148, 31, 220, 31, 31, 31, 103, 31, 144, 31, 178, 31, 236, 31, 236, 30, 236, 29, 236, 28, 236, 27, 236, 26, 236, 25, 236, 24, 236, 23, 236, 22, 236, 21, 236, 20, 236, 19, 236, 18, 236, 17, 236, 16, 236, 15, 236, 14, 236, 13, 236, 12, 236, 11, 236, 10, 236, 9, 236, 8, 236, 7, 236, 6, 236, 5, 236, 4, 236, 3, 236, 2, 162, 31, 121, 31, 199, 31, 149, 31, 167, 31, 45, 31, 254, 31, 154, 31, 163, 31, 146, 31, 34, 31, 190, 31, 155, 31, 241, 31, 143, 31, 34, 31, 165, 31, 58, 31, 17, 31, 44, 31, 63, 31, 70, 31, 164, 31, 47, 31, 3, 31, 236, 31, 177, 31, 158, 31, 220, 31, 179, 31, 1, 31, 240, 31, 218, 31, 139, 31, 149, 31, 166, 31, 243, 31, 208, 31, 123, 31, 140, 31, 8, 31, 66, 31, 51, 31, 162, 31, 135, 31, 19, 31, 143, 31, 172, 31, 248, 31, 16, 31, 77, 31, 103, 31, 102, 31, 78, 31, 78, 30, 78, 29, 78, 28, 78, 27, 78, 26, 78, 25, 78, 24, 78, 23, 78, 22, 78, 21, 78, 20, 78, 19, 78, 18, 78, 17, 78, 16, 78, 15, 78, 14, 78, 13, 78, 12, 78, 11, 78, 10, 78, 9, 78, 8, 78, 7, 78, 6, 78, 5, 78, 4, 78, 3, 78, 2, 78, 1, 78, 0, 78, 0, 78, 0, 78, 0, 78, 0, 219, 31, 196, 31, 25, 31, 2, 31, 163, 31, 204, 31, 125, 31, 50, 31, 56, 31, 206, 31, 70, 31, 32, 31, 32, 31, 61, 31, 158, 31, 56, 31, 166, 31, 223, 31, 111, 31, 95, 31, 83, 31, 225, 31, 229, 31, 84, 31, 134, 31, 94, 31, 9, 31, 53, 31, 129, 31, 119, 31, 118, 31, 244, 31, 250, 31, 159, 31, 190, 31, 200, 31, 115, 31, 134, 31, 72, 31, 205, 31, 105, 31, 154, 31, 168, 31, 133, 31, 109, 31, 185, 31, 54, 31, 36, 31, 121, 31, 26, 31, 74, 31, 4, 31, 13, 31, 250, 31, 77, 31, 151, 31, 28, 31, 113, 31, 194, 31, 56, 31, 81, 31, 51, 31, 131, 31, 21, 31, 162, 31, 121, 31, 125, 31, 212, 31, 255, 31, 123, 31, 163, 31, 102, 31, 253, 31, 76, 31, 201, 31, 233, 31, 232, 31, 178, 31, 178, 30, 178, 29, 178, 28, 178, 27, 178, 26, 178, 25, 178, 24, 178, 23, 178, 22, 178, 21, 178, 20, 178, 19, 178, 18, 178, 17, 178, 16, 178, 15, 178, 14, 78, 31, 87, 31, 44, 31, 220, 31, 157, 31, 81, 31, 180, 31, 174, 31, 38, 31, 89, 31, 234, 31, 109, 31, 122, 31, 3, 31, 41, 31, 214, 31, 162, 31, 123, 31, 94, 31, 220, 31, 107, 31, 1, 31, 26, 31, 187, 31, 97, 31, 13, 31, 238, 31, 163, 31, 6, 31, 119, 31, 31, 31, 20, 31, 161, 31, 218, 31, 130, 31, 43, 31, 254, 31, 145, 31, 247, 31, 6, 31, 200, 31, 30, 31, 13, 31, 81, 31, 101, 31, 205, 31, 12, 31, 201, 31, 255, 31, 11, 31, 234, 31, 90, 31, 201, 31, 253, 31, 211, 31, 72, 31, 23, 31, 98, 31, 23, 31, 182, 31, 243, 31, 74, 31, 239, 31, 239, 31, 147, 31, 180, 31, 140, 31, 239, 31, 66, 31, 181, 31, 42, 31, 219, 31, 24, 31, 70, 31, 234, 31, 92, 31, 145, 31, 143, 31, 143, 30, 143, 29, 143, 28, 143, 27, 143, 26, 143, 25, 143, 24, 143, 23, 143, 22, 143, 21, 143, 20, 143, 19, 143, 18, 143, 17, 143, 16, 143, 15, 143, 14, 143, 13, 143, 12, 143, 11, 143, 10, 143, 9, 143, 8, 143, 7, 143, 6, 143, 5, 143, 4, 143, 3, 143, 2, 143, 1, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 143, 0, 212, 31, 212, 30, 212, 29, 212, 28, 212, 27, 212, 26, 212, 25, 212, 24, 212, 23, 212, 22, 212, 21, 212, 20, 212, 19, 212, 18, 212, 17, 212, 16, 212, 15, 212, 14, 212, 13, 212, 12, 212, 11, 212, 10, 212, 9, 212, 8, 212, 7, 212, 6, 212, 5, 212, 4, 212, 3, 105, 31, 251, 31, 85, 31, 88, 31, 23, 31, 50, 31, 112, 31, 63, 31, 42, 31, 116, 31, 142, 31, 214, 31, 66, 31, 52, 31, 141, 31, 191, 31, 82, 31, 40, 31, 178, 31, 161, 31, 91, 31, 218, 31, 159, 31, 92, 31, 93, 31, 179, 31, 111, 31, 102, 31, 116, 31, 29, 31, 63, 31, 96, 31, 200, 31, 49, 31, 58, 31, 182, 31, 37, 31, 93, 31, 134, 31, 6, 31, 172, 31, 124, 31, 191, 31, 117, 31, 143, 31, 172, 31, 249, 31, 30, 31, 69, 31, 203, 31, 203, 30, 203, 29, 203, 28, 203, 27, 203, 26, 203, 25, 133, 31, 202, 31, 92, 31, 23, 31, 23, 31, 226, 31, 26, 31, 215, 31, 12, 31, 235, 31, 102, 31, 205, 31, 146, 31, 141, 31, 48, 31, 156, 31, 169, 31, 16, 31, 130, 31, 138, 31, 62, 31, 146, 31, 185, 31, 1, 31, 181, 31, 8, 31, 121, 31, 156, 31, 5, 31, 80, 31, 167, 31, 255, 31, 134, 31, 57, 31, 66, 31, 247, 31, 48, 31, 213, 31, 9, 31, 55, 31, 55, 31, 6, 31, 235, 31, 230, 31, 18, 31, 31, 31, 62, 31, 145, 31, 107, 31, 129, 31, 167, 31, 206, 31, 143, 31, 222, 31, 125, 31, 123, 31, 157, 31, 155, 31, 199, 31, 49, 31, 141, 31, 255, 31, 26, 31, 35, 31, 37, 31, 244, 31, 35, 31, 115, 31, 122, 31, 122, 30, 122, 29, 122, 28, 122, 27, 122, 26, 122, 25, 122, 24, 122, 23, 122, 22, 122, 21, 122, 20, 122, 19, 122, 18, 122, 17, 122, 16, 122, 15, 122, 14, 122, 13, 122, 12, 122, 11, 122, 10, 122, 9, 122, 8, 122, 7, 122, 6, 122, 5, 122, 4, 122, 3, 122, 2, 122, 1, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 122, 0, 208, 31, 74, 31, 116, 31, 177, 31, 228, 31, 44, 31, 200, 31, 255, 31, 134, 31, 108, 31, 35, 31, 194, 31, 223, 31, 119, 31, 105, 31, 30, 31, 35, 31, 196, 31, 157, 31, 109, 31, 209, 31, 204, 31, 204, 30, 79, 31, 17, 31, 201, 31, 253, 31, 46, 31, 131, 31, 131, 31, 252, 31, 122, 31, 200, 31, 159, 31, 193, 31, 10, 31, 196, 31, 139, 31, 224, 31, 210, 31, 2, 31, 212, 31, 153, 31, 32, 31, 225, 31, 33, 31, 8, 31, 5, 31, 245, 31, 152, 31, 132, 31, 28, 31, 66, 31, 60, 31, 213, 31, 127, 31, 14, 31, 101, 31, 172, 31, 124, 31, 91, 31, 154, 31, 194, 31, 193, 31, 22, 31, 127, 31, 110, 31, 49, 31, 179, 31, 22, 31, 135, 31, 119, 31, 141, 31, 97, 31, 64, 31, 23, 31, 56, 31, 144, 31, 221, 31, 12, 31, 244, 31, 61, 31, 65, 31, 156, 31, 102, 31, 228, 31, 195, 31, 35, 31, 32, 31, 206, 31, 57, 31, 129, 31, 148, 31, 38, 31, 89, 31, 89, 31, 239, 31, 191, 31, 165, 31, 73, 31, 64, 31, 128, 31, 155, 31, 41, 31, 217, 31, 195, 31, 221, 31, 31, 31, 181, 31, 160, 31, 161, 31, 41, 31, 144, 31, 128, 31, 236, 31, 46, 31, 163, 31, 69, 31, 50, 31, 9, 31, 171, 31, 239, 31, 186, 31, 57, 31, 192, 31, 197, 31, 176, 31, 2, 31, 157, 31, 200, 31, 90, 31, 76, 31, 52, 31);
    constant SCENARIO_ADDRESS_5 : integer := 40089;


    -- sixth run

    constant SCENARIO_LENGTH_K : integer := 0;
    constant SCENARIO_LENGTH_6 : integer := 1;
    type scenario_type_6 is array (0 to SCENARIO_LENGTH_6*2-1) of integer;
    signal scenario_input_6 : scenario_type_6 := (12, 13);
    signal scenario_full_6  : scenario_type_6 := (12, 13);
    constant SCENARIO_ADDRESS_6 : integer := 42089;


    -- seventh run

    constant SCENARIO_LENGTH_7 : integer := 1;
    type scenario_type_7 is array (0 to SCENARIO_LENGTH_7*2-1) of integer;
    signal scenario_input_7 : scenario_type_7 := (1, 1);
    signal scenario_full_7  : scenario_type_7 := (1, 1);
    constant SCENARIO_ADDRESS_7 : integer := 43089;



    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;


        -- Configure second run
        
        for i in 0 to SCENARIO_LENGTH_2*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_2+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_2(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        -- Configure third run

        for i in 0 to SCENARIO_LENGTH_3*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_3+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_3(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        -- Configure fourth run

        for i in 0 to SCENARIO_LENGTH_4*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_4+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_4(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        -- Configure fifth run

        for i in 0 to SCENARIO_LENGTH_5*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_5+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_5(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

         -- Configure sixth run

        for i in 0 to SCENARIO_LENGTH_6*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_6+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_6(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        -- Configure seventh run

        for i in 0 to SCENARIO_LENGTH_7*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_7+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_7(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;


        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';

        -- start sencond run without reset

        wait for 50 ns;

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_2, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_2, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';

        -- start third run without reset

        wait for 50 ns;

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_3, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_3, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
        
        wait for 5 ns;
        
        tb_start <= '0';


        -- start fourth run without reset

        wait for 100 ns;

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_4, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_4, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 90 ns;
        
        tb_start <= '0';


        -- start fifth run without reset

        wait for 100 ns;

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_5, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_5, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';


        -- start sixth run without reset

        wait for 50 ns;

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_6, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_K, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 100 ns;
        
        tb_start <= '0';


        -- start seventh run without reset

        wait for 50 ns;

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_7, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_K, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';

        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);


        -- second run
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH_2*2-1 loop
            assert RAM(SCENARIO_ADDRESS_2+i) = std_logic_vector(to_unsigned(scenario_full_2(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_2(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);



        -- third run
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH_3*2-1 loop
            assert RAM(SCENARIO_ADDRESS_3+i) = std_logic_vector(to_unsigned(scenario_full_3(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_3(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);


        -- fourth run
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH_4*2-1 loop
            assert RAM(SCENARIO_ADDRESS_4+i) = std_logic_vector(to_unsigned(scenario_full_4(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_4(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);


        -- fifth run
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH_5*2-1 loop
            assert RAM(SCENARIO_ADDRESS_5+i) = std_logic_vector(to_unsigned(scenario_full_5(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_5(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        -- sixth run
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH_6*2-1 loop
            assert RAM(SCENARIO_ADDRESS_6+i) = std_logic_vector(to_unsigned(scenario_full_6(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_6(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);


        -- seventh run
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH_7*2-1 loop
            assert RAM(SCENARIO_ADDRESS_7+i) = std_logic_vector(to_unsigned(scenario_full_7(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_7(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);



        -- end

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;
end architecture;
