-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_09 is
end project_tb_09;

architecture project_tb_09_arch of project_tb_09 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    signal memory_control : std_logic := '0';

    -- first run
    constant SCENARIO_LENGTH : integer := 737;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;
    signal scenario_input : scenario_type := (184, 0, 48, 0, 8, 0, 54, 0, 116, 0, 142, 0, 214, 0, 73, 0, 236, 0, 149, 0, 210, 0, 205, 0, 108, 0, 204, 0, 7, 0, 30, 0, 161, 0, 53, 0, 101, 0, 4, 0, 121, 0, 221, 0, 69, 0, 230, 0, 222, 0, 120, 0, 212, 0, 185, 0, 154, 0, 107, 0, 99, 0, 75, 0, 70, 0, 33, 0, 149, 0, 62, 0, 116, 0, 211, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 237, 0, 113, 0, 129, 0, 187, 0, 35, 0, 54, 0, 229, 0, 39, 0, 33, 0, 33, 0, 188, 0, 165, 0, 13, 0, 2, 0, 224, 0, 16, 0, 198, 0, 51, 0, 139, 0, 205, 0, 203, 0, 54, 0, 25, 0, 223, 0, 55, 0, 247, 0, 75, 0, 153, 0, 136, 0, 179, 0, 10, 0, 158, 0, 178, 0, 77, 0, 35, 0, 161, 0, 171, 0, 155, 0, 54, 0, 233, 0, 159, 0, 37, 0, 185, 0, 237, 0, 15, 0, 147, 0, 210, 0, 136, 0, 5, 0, 12, 0, 4, 0, 0, 0, 233, 0, 194, 0, 253, 0, 117, 0, 230, 0, 208, 0, 60, 0, 168, 0, 159, 0, 117, 0, 223, 0, 122, 0, 101, 0, 58, 0, 129, 0, 98, 0, 234, 0, 157, 0, 15, 0, 99, 0, 38, 0, 134, 0, 39, 0, 32, 0, 208, 0, 215, 0, 5, 0, 156, 0, 105, 0, 63, 0, 50, 0, 143, 0, 150, 0, 189, 0, 210, 0, 7, 0, 248, 0, 236, 0, 29, 0, 28, 0, 176, 0, 244, 0, 13, 0, 135, 0, 248, 0, 106, 0, 202, 0, 197, 0, 117, 0, 14, 0, 108, 0, 253, 0, 217, 0, 205, 0, 237, 0, 78, 0, 246, 0, 126, 0, 77, 0, 255, 0, 165, 0, 229, 0, 197, 0, 41, 0, 24, 0, 28, 0, 23, 0, 70, 0, 45, 0, 33, 0, 103, 0, 29, 0, 94, 0, 70, 0, 44, 0, 67, 0, 221, 0, 170, 0, 228, 0, 72, 0, 205, 0, 222, 0, 6, 0, 180, 0, 130, 0, 10, 0, 214, 0, 148, 0, 68, 0, 231, 0, 26, 0, 141, 0, 138, 0, 148, 0, 225, 0, 15, 0, 27, 0, 65, 0, 254, 0, 57, 0, 87, 0, 51, 0, 231, 0, 167, 0, 246, 0, 124, 0, 91, 0, 218, 0, 8, 0, 125, 0, 16, 0, 100, 0, 121, 0, 114, 0, 9, 0, 142, 0, 200, 0, 80, 0, 104, 0, 160, 0, 118, 0, 228, 0, 235, 0, 91, 0, 48, 0, 28, 0, 131, 0, 222, 0, 208, 0, 9, 0, 14, 0, 71, 0, 222, 0, 217, 0, 217, 0, 156, 0, 26, 0, 168, 0, 240, 0, 110, 0, 159, 0, 230, 0, 130, 0, 187, 0, 98, 0, 93, 0, 32, 0, 89, 0, 111, 0, 245, 0, 11, 0, 124, 0, 160, 0, 216, 0, 87, 0, 201, 0, 78, 0, 245, 0, 212, 0, 31, 0, 218, 0, 104, 0, 140, 0, 196, 0, 159, 0, 70, 0, 145, 0, 216, 0, 141, 0, 3, 0, 20, 0, 227, 0, 49, 0, 163, 0, 98, 0, 12, 0, 206, 0, 223, 0, 166, 0, 69, 0, 21, 0, 179, 0, 53, 0, 38, 0, 243, 0, 224, 0, 185, 0, 152, 0, 16, 0, 64, 0, 138, 0, 107, 0, 219, 0, 167, 0, 63, 0, 162, 0, 138, 0, 15, 0, 23, 0, 150, 0, 242, 0, 159, 0, 140, 0, 250, 0, 72, 0, 98, 0, 124, 0, 238, 0, 223, 0, 56, 0, 188, 0, 164, 0, 80, 0, 155, 0, 138, 0, 229, 0, 58, 0, 175, 0, 157, 0, 216, 0, 61, 0, 122, 0, 210, 0, 88, 0, 123, 0, 129, 0, 144, 0, 95, 0, 79, 0, 112, 0, 112, 0, 208, 0, 13, 0, 69, 0, 194, 0, 16, 0, 2, 0, 58, 0, 60, 0, 146, 0, 160, 0, 47, 0, 11, 0, 137, 0, 167, 0, 58, 0, 14, 0, 43, 0, 27, 0, 191, 0, 207, 0, 54, 0, 177, 0, 135, 0, 229, 0, 142, 0, 245, 0, 87, 0, 142, 0, 38, 0, 72, 0, 111, 0, 9, 0, 189, 0, 8, 0, 221, 0, 111, 0, 174, 0, 89, 0, 202, 0, 8, 0, 104, 0, 205, 0, 53, 0, 21, 0, 34, 0, 149, 0, 146, 0, 80, 0, 181, 0, 145, 0, 9, 0, 198, 0, 215, 0, 176, 0, 165, 0, 148, 0, 86, 0, 255, 0, 158, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 181, 0, 99, 0, 81, 0, 234, 0, 54, 0, 132, 0, 253, 0, 147, 0, 217, 0, 137, 0, 157, 0, 200, 0, 153, 0, 109, 0, 45, 0, 239, 0, 187, 0, 172, 0, 9, 0, 197, 0, 102, 0, 221, 0, 159, 0, 13, 0, 111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 0, 165, 0, 160, 0, 179, 0, 135, 0, 107, 0, 239, 0, 156, 0, 207, 0, 212, 0, 61, 0, 233, 0, 53, 0, 247, 0, 35, 0, 242, 0, 64, 0, 212, 0, 62, 0, 210, 0, 221, 0, 98, 0, 141, 0, 53, 0, 219, 0, 206, 0, 25, 0, 92, 0, 120, 0, 11, 0, 3, 0, 214, 0, 243, 0, 108, 0, 130, 0, 137, 0, 190, 0, 152, 0, 74, 0, 59, 0, 207, 0, 98, 0, 41, 0, 146, 0, 126, 0, 70, 0, 99, 0, 200, 0, 12, 0, 218, 0, 139, 0, 149, 0, 234, 0, 183, 0, 9, 0, 63, 0, 24, 0, 54, 0, 107, 0, 43, 0, 173, 0, 121, 0, 250, 0, 240, 0, 57, 0, 44, 0, 220, 0, 255, 0, 124, 0, 131, 0, 140, 0, 251, 0, 213, 0, 37, 0, 218, 0, 153, 0, 229, 0, 194, 0, 36, 0, 172, 0, 34, 0, 214, 0, 111, 0, 213, 0, 244, 0, 100, 0, 88, 0, 196, 0, 155, 0, 243, 0, 56, 0, 36, 0, 52, 0, 94, 0, 56, 0, 81, 0, 127, 0, 163, 0, 198, 0, 172, 0, 165, 0, 66, 0, 44, 0, 193, 0, 53, 0, 249, 0, 2, 0, 64, 0, 227, 0, 131, 0, 86, 0, 43, 0, 247, 0, 121, 0, 206, 0, 34, 0, 167, 0, 86, 0, 68, 0, 77, 0, 131, 0, 255, 0, 251, 0, 82, 0, 169, 0, 229, 0, 33, 0, 32, 0, 152, 0, 49, 0, 155, 0, 227, 0, 143, 0, 83, 0, 150, 0, 25, 0, 39, 0, 143, 0, 223, 0, 57, 0, 220, 0, 63, 0, 137, 0, 221, 0, 109, 0, 128, 0, 54, 0, 146, 0, 207, 0, 142, 0, 247, 0, 63, 0, 4, 0, 98, 0, 133, 0, 127, 0, 222, 0, 237, 0, 137, 0, 214, 0, 255, 0, 164, 0, 27, 0, 115, 0, 203, 0, 228, 0, 153, 0, 81, 0, 17, 0, 212, 0, 179, 0, 116, 0, 242, 0, 207, 0, 32, 0, 119, 0, 74, 0, 164, 0, 143, 0, 249, 0, 23, 0, 35, 0, 164, 0, 182, 0, 211, 0, 49, 0, 90, 0, 21, 0, 246, 0, 239, 0, 156, 0, 156, 0, 112, 0, 55, 0, 246, 0, 77, 0, 44, 0, 71, 0, 111, 0, 67, 0, 17, 0, 221, 0);
    signal scenario_full  : scenario_type := (184, 31, 48, 31, 8, 31, 54, 31, 116, 31, 142, 31, 214, 31, 73, 31, 236, 31, 149, 31, 210, 31, 205, 31, 108, 31, 204, 31, 7, 31, 30, 31, 161, 31, 53, 31, 101, 31, 4, 31, 121, 31, 221, 31, 69, 31, 230, 31, 222, 31, 120, 31, 212, 31, 185, 31, 154, 31, 107, 31, 99, 31, 75, 31, 70, 31, 33, 31, 149, 31, 62, 31, 116, 31, 211, 31, 211, 30, 211, 29, 211, 28, 211, 27, 211, 26, 211, 25, 211, 24, 211, 23, 211, 22, 211, 21, 211, 20, 211, 19, 211, 18, 211, 17, 211, 16, 211, 15, 211, 14, 211, 13, 211, 12, 211, 11, 211, 10, 211, 9, 211, 8, 211, 7, 211, 6, 211, 5, 211, 4, 211, 3, 211, 2, 211, 1, 237, 31, 113, 31, 129, 31, 187, 31, 35, 31, 54, 31, 229, 31, 39, 31, 33, 31, 33, 31, 188, 31, 165, 31, 13, 31, 2, 31, 224, 31, 16, 31, 198, 31, 51, 31, 139, 31, 205, 31, 203, 31, 54, 31, 25, 31, 223, 31, 55, 31, 247, 31, 75, 31, 153, 31, 136, 31, 179, 31, 10, 31, 158, 31, 178, 31, 77, 31, 35, 31, 161, 31, 171, 31, 155, 31, 54, 31, 233, 31, 159, 31, 37, 31, 185, 31, 237, 31, 15, 31, 147, 31, 210, 31, 136, 31, 5, 31, 12, 31, 4, 31, 4, 30, 233, 31, 194, 31, 253, 31, 117, 31, 230, 31, 208, 31, 60, 31, 168, 31, 159, 31, 117, 31, 223, 31, 122, 31, 101, 31, 58, 31, 129, 31, 98, 31, 234, 31, 157, 31, 15, 31, 99, 31, 38, 31, 134, 31, 39, 31, 32, 31, 208, 31, 215, 31, 5, 31, 156, 31, 105, 31, 63, 31, 50, 31, 143, 31, 150, 31, 189, 31, 210, 31, 7, 31, 248, 31, 236, 31, 29, 31, 28, 31, 176, 31, 244, 31, 13, 31, 135, 31, 248, 31, 106, 31, 202, 31, 197, 31, 117, 31, 14, 31, 108, 31, 253, 31, 217, 31, 205, 31, 237, 31, 78, 31, 246, 31, 126, 31, 77, 31, 255, 31, 165, 31, 229, 31, 197, 31, 41, 31, 24, 31, 28, 31, 23, 31, 70, 31, 45, 31, 33, 31, 103, 31, 29, 31, 94, 31, 70, 31, 44, 31, 67, 31, 221, 31, 170, 31, 228, 31, 72, 31, 205, 31, 222, 31, 6, 31, 180, 31, 130, 31, 10, 31, 214, 31, 148, 31, 68, 31, 231, 31, 26, 31, 141, 31, 138, 31, 148, 31, 225, 31, 15, 31, 27, 31, 65, 31, 254, 31, 57, 31, 87, 31, 51, 31, 231, 31, 167, 31, 246, 31, 124, 31, 91, 31, 218, 31, 8, 31, 125, 31, 16, 31, 100, 31, 121, 31, 114, 31, 9, 31, 142, 31, 200, 31, 80, 31, 104, 31, 160, 31, 118, 31, 228, 31, 235, 31, 91, 31, 48, 31, 28, 31, 131, 31, 222, 31, 208, 31, 9, 31, 14, 31, 71, 31, 222, 31, 217, 31, 217, 31, 156, 31, 26, 31, 168, 31, 240, 31, 110, 31, 159, 31, 230, 31, 130, 31, 187, 31, 98, 31, 93, 31, 32, 31, 89, 31, 111, 31, 245, 31, 11, 31, 124, 31, 160, 31, 216, 31, 87, 31, 201, 31, 78, 31, 245, 31, 212, 31, 31, 31, 218, 31, 104, 31, 140, 31, 196, 31, 159, 31, 70, 31, 145, 31, 216, 31, 141, 31, 3, 31, 20, 31, 227, 31, 49, 31, 163, 31, 98, 31, 12, 31, 206, 31, 223, 31, 166, 31, 69, 31, 21, 31, 179, 31, 53, 31, 38, 31, 243, 31, 224, 31, 185, 31, 152, 31, 16, 31, 64, 31, 138, 31, 107, 31, 219, 31, 167, 31, 63, 31, 162, 31, 138, 31, 15, 31, 23, 31, 150, 31, 242, 31, 159, 31, 140, 31, 250, 31, 72, 31, 98, 31, 124, 31, 238, 31, 223, 31, 56, 31, 188, 31, 164, 31, 80, 31, 155, 31, 138, 31, 229, 31, 58, 31, 175, 31, 157, 31, 216, 31, 61, 31, 122, 31, 210, 31, 88, 31, 123, 31, 129, 31, 144, 31, 95, 31, 79, 31, 112, 31, 112, 31, 208, 31, 13, 31, 69, 31, 194, 31, 16, 31, 2, 31, 58, 31, 60, 31, 146, 31, 160, 31, 47, 31, 11, 31, 137, 31, 167, 31, 58, 31, 14, 31, 43, 31, 27, 31, 191, 31, 207, 31, 54, 31, 177, 31, 135, 31, 229, 31, 142, 31, 245, 31, 87, 31, 142, 31, 38, 31, 72, 31, 111, 31, 9, 31, 189, 31, 8, 31, 221, 31, 111, 31, 174, 31, 89, 31, 202, 31, 8, 31, 104, 31, 205, 31, 53, 31, 21, 31, 34, 31, 149, 31, 146, 31, 80, 31, 181, 31, 145, 31, 9, 31, 198, 31, 215, 31, 176, 31, 165, 31, 148, 31, 86, 31, 255, 31, 158, 31, 158, 30, 158, 29, 158, 28, 158, 27, 158, 26, 158, 25, 158, 24, 158, 23, 158, 22, 158, 21, 158, 20, 158, 19, 158, 18, 158, 17, 158, 16, 158, 15, 158, 14, 158, 13, 158, 12, 158, 11, 158, 10, 158, 9, 158, 8, 158, 7, 158, 6, 158, 5, 158, 4, 158, 3, 158, 2, 158, 1, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 158, 0, 181, 31, 99, 31, 81, 31, 234, 31, 54, 31, 132, 31, 253, 31, 147, 31, 217, 31, 137, 31, 157, 31, 200, 31, 153, 31, 109, 31, 45, 31, 239, 31, 187, 31, 172, 31, 9, 31, 197, 31, 102, 31, 221, 31, 159, 31, 13, 31, 111, 31, 111, 30, 111, 29, 111, 28, 111, 27, 111, 26, 111, 25, 111, 24, 111, 23, 111, 22, 111, 21, 111, 20, 111, 19, 111, 18, 111, 17, 111, 16, 111, 15, 111, 14, 111, 13, 111, 12, 111, 11, 111, 10, 111, 9, 111, 8, 111, 7, 111, 6, 111, 5, 111, 4, 111, 3, 111, 2, 111, 1, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 111, 0, 66, 31, 165, 31, 160, 31, 179, 31, 135, 31, 107, 31, 239, 31, 156, 31, 207, 31, 212, 31, 61, 31, 233, 31, 53, 31, 247, 31, 35, 31, 242, 31, 64, 31, 212, 31, 62, 31, 210, 31, 221, 31, 98, 31, 141, 31, 53, 31, 219, 31, 206, 31, 25, 31, 92, 31, 120, 31, 11, 31, 3, 31, 214, 31, 243, 31, 108, 31, 130, 31, 137, 31, 190, 31, 152, 31, 74, 31, 59, 31, 207, 31, 98, 31, 41, 31, 146, 31, 126, 31, 70, 31, 99, 31, 200, 31, 12, 31, 218, 31, 139, 31, 149, 31, 234, 31, 183, 31, 9, 31, 63, 31, 24, 31, 54, 31, 107, 31, 43, 31, 173, 31, 121, 31, 250, 31, 240, 31, 57, 31, 44, 31, 220, 31, 255, 31, 124, 31, 131, 31, 140, 31, 251, 31, 213, 31, 37, 31, 218, 31, 153, 31, 229, 31, 194, 31, 36, 31, 172, 31, 34, 31, 214, 31, 111, 31, 213, 31, 244, 31, 100, 31, 88, 31, 196, 31, 155, 31, 243, 31, 56, 31, 36, 31, 52, 31, 94, 31, 56, 31, 81, 31, 127, 31, 163, 31, 198, 31, 172, 31, 165, 31, 66, 31, 44, 31, 193, 31, 53, 31, 249, 31, 2, 31, 64, 31, 227, 31, 131, 31, 86, 31, 43, 31, 247, 31, 121, 31, 206, 31, 34, 31, 167, 31, 86, 31, 68, 31, 77, 31, 131, 31, 255, 31, 251, 31, 82, 31, 169, 31, 229, 31, 33, 31, 32, 31, 152, 31, 49, 31, 155, 31, 227, 31, 143, 31, 83, 31, 150, 31, 25, 31, 39, 31, 143, 31, 223, 31, 57, 31, 220, 31, 63, 31, 137, 31, 221, 31, 109, 31, 128, 31, 54, 31, 146, 31, 207, 31, 142, 31, 247, 31, 63, 31, 4, 31, 98, 31, 133, 31, 127, 31, 222, 31, 237, 31, 137, 31, 214, 31, 255, 31, 164, 31, 27, 31, 115, 31, 203, 31, 228, 31, 153, 31, 81, 31, 17, 31, 212, 31, 179, 31, 116, 31, 242, 31, 207, 31, 32, 31, 119, 31, 74, 31, 164, 31, 143, 31, 249, 31, 23, 31, 35, 31, 164, 31, 182, 31, 211, 31, 49, 31, 90, 31, 21, 31, 246, 31, 239, 31, 156, 31, 156, 31, 112, 31, 55, 31, 246, 31, 77, 31, 44, 31, 71, 31, 111, 31, 67, 31, 17, 31, 221, 31);
    constant SCENARIO_ADDRESS : integer := 890;

    -- second run

    constant SCENARIO_LENGTH_2 : integer := 1022;
    type scenario_type_2 is array (0 to SCENARIO_LENGTH_2*2-1) of integer;
    signal scenario_input_2 : scenario_type_2 := (102, 0, 192, 0, 194, 0, 31, 0, 186, 0, 142, 0, 159, 0, 46, 0, 140, 0, 108, 0, 53, 0, 29, 0, 172, 0, 87, 0, 9, 0, 56, 0, 6, 0, 229, 0, 163, 0, 85, 0, 195, 0, 30, 0, 203, 0, 117, 0, 152, 0, 164, 0, 82, 0, 144, 0, 128, 0, 76, 0, 56, 0, 248, 0, 66, 0, 95, 0, 240, 0, 201, 0, 197, 0, 204, 0, 223, 0, 40, 0, 208, 0, 4, 0, 71, 0, 113, 0, 79, 0, 243, 0, 145, 0, 212, 0, 40, 0, 160, 0, 202, 0, 80, 0, 230, 0, 117, 0, 37, 0, 190, 0, 199, 0, 82, 0, 29, 0, 191, 0, 155, 0, 24, 0, 144, 0, 124, 0, 124, 0, 91, 0, 173, 0, 95, 0, 233, 0, 69, 0, 137, 0, 24, 0, 51, 0, 238, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 191, 0, 110, 0, 118, 0, 13, 0, 198, 0, 100, 0, 53, 0, 160, 0, 127, 0, 195, 0, 119, 0, 166, 0, 29, 0, 61, 0, 52, 0, 68, 0, 129, 0, 174, 0, 221, 0, 157, 0, 232, 0, 43, 0, 103, 0, 140, 0, 104, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 142, 0, 107, 0, 99, 0, 166, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 229, 0, 66, 0, 115, 0, 175, 0, 68, 0, 29, 0, 252, 0, 77, 0, 147, 0, 245, 0, 157, 0, 16, 0, 28, 0, 243, 0, 236, 0, 223, 0, 16, 0, 39, 0, 212, 0, 206, 0, 183, 0, 64, 0, 78, 0, 195, 0, 158, 0, 60, 0, 14, 0, 183, 0, 206, 0, 121, 0, 126, 0, 160, 0, 49, 0, 120, 0, 60, 0, 63, 0, 204, 0, 152, 0, 110, 0, 122, 0, 193, 0, 214, 0, 2, 0, 226, 0, 102, 0, 88, 0, 243, 0, 10, 0, 191, 0, 180, 0, 11, 0, 236, 0, 181, 0, 73, 0, 138, 0, 75, 0, 172, 0, 62, 0, 58, 0, 107, 0, 46, 0, 90, 0, 215, 0, 4, 0, 227, 0, 29, 0, 161, 0, 43, 0, 2, 0, 19, 0, 86, 0, 174, 0, 195, 0, 106, 0, 144, 0, 29, 0, 87, 0, 219, 0, 60, 0, 170, 0, 171, 0, 148, 0, 22, 0, 53, 0, 76, 0, 142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 252, 0, 54, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 139, 0, 99, 0, 221, 0, 162, 0, 151, 0, 164, 0, 96, 0, 32, 0, 128, 0, 118, 0, 168, 0, 200, 0, 97, 0, 57, 0, 145, 0, 84, 0, 74, 0, 125, 0, 164, 0, 10, 0, 203, 0, 8, 0, 68, 0, 247, 0, 12, 0, 220, 0, 95, 0, 22, 0, 213, 0, 67, 0, 60, 0, 196, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 163, 0, 233, 0, 66, 0, 82, 0, 102, 0, 196, 0, 214, 0, 134, 0, 196, 0, 180, 0, 24, 0, 250, 0, 27, 0, 92, 0, 200, 0, 239, 0, 243, 0, 175, 0, 80, 0, 43, 0, 19, 0, 176, 0, 119, 0, 168, 0, 247, 0, 117, 0, 253, 0, 240, 0, 51, 0, 115, 0, 188, 0, 222, 0, 101, 0, 207, 0, 84, 0, 7, 0, 252, 0, 177, 0, 171, 0, 175, 0, 222, 0, 209, 0, 188, 0, 199, 0, 116, 0, 39, 0, 49, 0, 230, 0, 184, 0, 112, 0, 200, 0, 203, 0, 45, 0, 134, 0, 3, 0, 20, 0, 245, 0, 68, 0, 238, 0, 76, 0, 125, 0, 93, 0, 150, 0, 103, 0, 185, 0, 89, 0, 166, 0, 159, 0, 33, 0, 235, 0, 247, 0, 187, 0, 57, 0, 247, 0, 249, 0, 104, 0, 201, 0, 251, 0, 51, 0, 102, 0, 73, 0, 223, 0, 75, 0, 242, 0, 137, 0, 139, 0, 161, 0, 189, 0, 178, 0, 247, 0, 85, 0, 131, 0, 181, 0, 250, 0, 138, 0, 47, 0, 139, 0, 67, 0, 62, 0, 32, 0, 62, 0, 178, 0, 62, 0, 75, 0, 197, 0, 122, 0, 72, 0, 25, 0, 60, 0, 208, 0, 0, 0, 186, 0, 133, 0, 190, 0, 154, 0, 179, 0, 233, 0, 112, 0, 40, 0, 15, 0, 251, 0, 112, 0, 233, 0, 233, 0, 195, 0, 247, 0, 152, 0, 43, 0, 204, 0, 44, 0, 145, 0, 81, 0, 163, 0, 162, 0, 102, 0, 220, 0, 77, 0, 96, 0, 219, 0, 12, 0, 136, 0, 3, 0, 134, 0, 95, 0, 85, 0, 26, 0, 176, 0, 129, 0, 164, 0, 160, 0, 252, 0, 66, 0, 148, 0, 51, 0, 208, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 100, 0, 2, 0, 131, 0, 242, 0, 77, 0, 192, 0, 85, 0, 166, 0, 105, 0, 126, 0, 10, 0, 53, 0, 93, 0, 193, 0, 162, 0, 79, 0, 160, 0, 221, 0, 214, 0, 235, 0, 69, 0, 147, 0, 222, 0, 93, 0, 44, 0, 208, 0, 133, 0, 94, 0, 177, 0, 104, 0, 111, 0, 203, 0, 58, 0, 105, 0, 9, 0, 176, 0, 1, 0, 164, 0, 123, 0, 33, 0, 219, 0, 165, 0, 175, 0, 21, 0, 18, 0, 182, 0, 136, 0, 246, 0, 15, 0, 232, 0, 12, 0, 233, 0, 20, 0, 46, 0, 20, 0, 180, 0, 61, 0, 207, 0, 23, 0, 100, 0, 129, 0, 249, 0, 156, 0, 200, 0, 173, 0, 64, 0, 233, 0, 133, 0, 169, 0, 94, 0, 121, 0, 13, 0, 77, 0, 84, 0, 200, 0, 121, 0, 70, 0, 50, 0, 254, 0, 19, 0, 228, 0, 53, 0, 158, 0, 47, 0, 250, 0, 220, 0, 238, 0, 161, 0, 218, 0, 73, 0, 145, 0, 54, 0, 248, 0, 89, 0, 40, 0, 27, 0, 235, 0, 177, 0, 233, 0, 43, 0, 12, 0, 174, 0, 135, 0, 8, 0, 171, 0, 100, 0, 54, 0, 195, 0, 250, 0, 96, 0, 25, 0, 189, 0, 155, 0, 102, 0, 229, 0, 37, 0, 212, 0, 113, 0, 196, 0, 137, 0, 202, 0, 73, 0, 157, 0, 242, 0, 176, 0, 87, 0, 164, 0, 186, 0, 52, 0, 240, 0, 69, 0, 10, 0, 100, 0, 39, 0, 90, 0, 138, 0, 110, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 186, 0, 246, 0, 254, 0, 127, 0, 195, 0, 71, 0, 197, 0, 235, 0, 125, 0, 8, 0, 2, 0, 201, 0, 94, 0, 228, 0, 124, 0, 230, 0, 56, 0, 111, 0, 158, 0, 48, 0, 132, 0, 144, 0, 6, 0, 128, 0, 171, 0, 200, 0, 187, 0, 80, 0, 68, 0, 54, 0, 125, 0, 104, 0, 131, 0, 126, 0, 224, 0, 178, 0, 54, 0, 143, 0, 206, 0, 16, 0, 227, 0, 164, 0, 38, 0, 41, 0, 165, 0, 55, 0, 251, 0, 73, 0, 169, 0, 187, 0, 198, 0, 194, 0, 72, 0, 183, 0, 123, 0, 240, 0, 198, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 150, 0, 44, 0, 35, 0, 226, 0, 29, 0, 100, 0, 128, 0, 76, 0, 198, 0, 201, 0, 121, 0, 99, 0, 116, 0, 203, 0, 144, 0, 18, 0, 248, 0, 203, 0, 6, 0, 132, 0, 124, 0, 139, 0, 22, 0, 28, 0, 0, 0, 173, 0, 215, 0, 64, 0, 201, 0, 184, 0, 90, 0, 69, 0, 60, 0, 81, 0, 18, 0, 38, 0, 167, 0, 79, 0, 28, 0, 222, 0, 85, 0, 69, 0, 239, 0, 73, 0, 224, 0, 38, 0, 179, 0, 198, 0, 244, 0, 62, 0, 227, 0, 193, 0, 30, 0, 28, 0, 68, 0, 15, 0, 4, 0, 128, 0, 79, 0, 247, 0, 54, 0, 215, 0, 39, 0, 198, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 121, 0, 168, 0, 105, 0, 73, 0, 53, 0, 210, 0, 71, 0, 157, 0, 229, 0, 98, 0, 117, 0, 247, 0, 241, 0, 43, 0, 156, 0, 139, 0, 81, 0, 46, 0, 54, 0, 129, 0, 90, 0, 27, 0, 250, 0, 247, 0, 146, 0, 202, 0, 119, 0, 227, 0, 5, 0, 67, 0, 145, 0, 237, 0, 12, 0, 144, 0, 40, 0, 153, 0, 223, 0, 129, 0, 155, 0, 26, 0, 233, 0, 255, 0, 205, 0, 79, 0, 48, 0, 168, 0, 63, 0, 73, 0, 154, 0, 130, 0, 162, 0, 64, 0, 84, 0, 72, 0, 124, 0, 73, 0, 155, 0, 33, 0, 51, 0, 209, 0, 119, 0, 204, 0, 58, 0, 41, 0);
    signal scenario_full_2  : scenario_type_2 := (102, 31, 192, 31, 194, 31, 31, 31, 186, 31, 142, 31, 159, 31, 46, 31, 140, 31, 108, 31, 53, 31, 29, 31, 172, 31, 87, 31, 9, 31, 56, 31, 6, 31, 229, 31, 163, 31, 85, 31, 195, 31, 30, 31, 203, 31, 117, 31, 152, 31, 164, 31, 82, 31, 144, 31, 128, 31, 76, 31, 56, 31, 248, 31, 66, 31, 95, 31, 240, 31, 201, 31, 197, 31, 204, 31, 223, 31, 40, 31, 208, 31, 4, 31, 71, 31, 113, 31, 79, 31, 243, 31, 145, 31, 212, 31, 40, 31, 160, 31, 202, 31, 80, 31, 230, 31, 117, 31, 37, 31, 190, 31, 199, 31, 82, 31, 29, 31, 191, 31, 155, 31, 24, 31, 144, 31, 124, 31, 124, 31, 91, 31, 173, 31, 95, 31, 233, 31, 69, 31, 137, 31, 24, 31, 51, 31, 238, 31, 238, 30, 238, 29, 238, 28, 238, 27, 238, 26, 238, 25, 238, 24, 238, 23, 238, 22, 238, 21, 238, 20, 238, 19, 238, 18, 238, 17, 238, 16, 238, 15, 238, 14, 238, 13, 238, 12, 238, 11, 238, 10, 238, 9, 238, 8, 238, 7, 238, 6, 238, 5, 238, 4, 238, 3, 238, 2, 238, 1, 238, 0, 238, 0, 238, 0, 238, 0, 238, 0, 238, 0, 238, 0, 238, 0, 238, 0, 238, 0, 238, 0, 238, 0, 191, 31, 110, 31, 118, 31, 13, 31, 198, 31, 100, 31, 53, 31, 160, 31, 127, 31, 195, 31, 119, 31, 166, 31, 29, 31, 61, 31, 52, 31, 68, 31, 129, 31, 174, 31, 221, 31, 157, 31, 232, 31, 43, 31, 103, 31, 140, 31, 104, 31, 104, 30, 104, 29, 104, 28, 104, 27, 104, 26, 104, 25, 104, 24, 104, 23, 104, 22, 104, 21, 104, 20, 104, 19, 104, 18, 104, 17, 104, 16, 104, 15, 104, 14, 104, 13, 104, 12, 104, 11, 104, 10, 104, 9, 104, 8, 104, 7, 104, 6, 104, 5, 104, 4, 104, 3, 104, 2, 104, 1, 104, 0, 104, 0, 104, 0, 142, 31, 107, 31, 99, 31, 166, 31, 25, 31, 25, 30, 25, 29, 25, 28, 25, 27, 25, 26, 25, 25, 25, 24, 25, 23, 25, 22, 25, 21, 25, 20, 25, 19, 25, 18, 25, 17, 25, 16, 25, 15, 25, 14, 25, 13, 25, 12, 25, 11, 25, 10, 25, 9, 25, 8, 25, 7, 25, 6, 25, 5, 25, 4, 25, 3, 25, 2, 25, 1, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 25, 0, 229, 31, 66, 31, 115, 31, 175, 31, 68, 31, 29, 31, 252, 31, 77, 31, 147, 31, 245, 31, 157, 31, 16, 31, 28, 31, 243, 31, 236, 31, 223, 31, 16, 31, 39, 31, 212, 31, 206, 31, 183, 31, 64, 31, 78, 31, 195, 31, 158, 31, 60, 31, 14, 31, 183, 31, 206, 31, 121, 31, 126, 31, 160, 31, 49, 31, 120, 31, 60, 31, 63, 31, 204, 31, 152, 31, 110, 31, 122, 31, 193, 31, 214, 31, 2, 31, 226, 31, 102, 31, 88, 31, 243, 31, 10, 31, 191, 31, 180, 31, 11, 31, 236, 31, 181, 31, 73, 31, 138, 31, 75, 31, 172, 31, 62, 31, 58, 31, 107, 31, 46, 31, 90, 31, 215, 31, 4, 31, 227, 31, 29, 31, 161, 31, 43, 31, 2, 31, 19, 31, 86, 31, 174, 31, 195, 31, 106, 31, 144, 31, 29, 31, 87, 31, 219, 31, 60, 31, 170, 31, 171, 31, 148, 31, 22, 31, 53, 31, 76, 31, 142, 31, 142, 30, 142, 29, 142, 28, 142, 27, 142, 26, 142, 25, 142, 24, 142, 23, 142, 22, 142, 21, 142, 20, 142, 19, 142, 18, 142, 17, 142, 16, 142, 15, 142, 14, 142, 13, 142, 12, 142, 11, 142, 10, 142, 9, 142, 8, 142, 7, 142, 6, 142, 5, 142, 4, 142, 3, 142, 2, 142, 1, 142, 0, 142, 0, 142, 0, 142, 0, 142, 0, 142, 0, 142, 0, 142, 0, 142, 0, 142, 0, 142, 0, 142, 0, 142, 0, 252, 31, 54, 31, 30, 31, 30, 30, 30, 29, 30, 28, 30, 27, 30, 26, 30, 25, 30, 24, 30, 23, 30, 22, 30, 21, 30, 20, 30, 19, 30, 18, 30, 17, 30, 16, 30, 15, 30, 14, 30, 13, 30, 12, 30, 11, 139, 31, 99, 31, 221, 31, 162, 31, 151, 31, 164, 31, 96, 31, 32, 31, 128, 31, 118, 31, 168, 31, 200, 31, 97, 31, 57, 31, 145, 31, 84, 31, 74, 31, 125, 31, 164, 31, 10, 31, 203, 31, 8, 31, 68, 31, 247, 31, 12, 31, 220, 31, 95, 31, 22, 31, 213, 31, 67, 31, 60, 31, 196, 31, 196, 30, 196, 29, 196, 28, 196, 27, 196, 26, 196, 25, 196, 24, 196, 23, 196, 22, 196, 21, 196, 20, 196, 19, 163, 31, 233, 31, 66, 31, 82, 31, 102, 31, 196, 31, 214, 31, 134, 31, 196, 31, 180, 31, 24, 31, 250, 31, 27, 31, 92, 31, 200, 31, 239, 31, 243, 31, 175, 31, 80, 31, 43, 31, 19, 31, 176, 31, 119, 31, 168, 31, 247, 31, 117, 31, 253, 31, 240, 31, 51, 31, 115, 31, 188, 31, 222, 31, 101, 31, 207, 31, 84, 31, 7, 31, 252, 31, 177, 31, 171, 31, 175, 31, 222, 31, 209, 31, 188, 31, 199, 31, 116, 31, 39, 31, 49, 31, 230, 31, 184, 31, 112, 31, 200, 31, 203, 31, 45, 31, 134, 31, 3, 31, 20, 31, 245, 31, 68, 31, 238, 31, 76, 31, 125, 31, 93, 31, 150, 31, 103, 31, 185, 31, 89, 31, 166, 31, 159, 31, 33, 31, 235, 31, 247, 31, 187, 31, 57, 31, 247, 31, 249, 31, 104, 31, 201, 31, 251, 31, 51, 31, 102, 31, 73, 31, 223, 31, 75, 31, 242, 31, 137, 31, 139, 31, 161, 31, 189, 31, 178, 31, 247, 31, 85, 31, 131, 31, 181, 31, 250, 31, 138, 31, 47, 31, 139, 31, 67, 31, 62, 31, 32, 31, 62, 31, 178, 31, 62, 31, 75, 31, 197, 31, 122, 31, 72, 31, 25, 31, 60, 31, 208, 31, 208, 30, 186, 31, 133, 31, 190, 31, 154, 31, 179, 31, 233, 31, 112, 31, 40, 31, 15, 31, 251, 31, 112, 31, 233, 31, 233, 31, 195, 31, 247, 31, 152, 31, 43, 31, 204, 31, 44, 31, 145, 31, 81, 31, 163, 31, 162, 31, 102, 31, 220, 31, 77, 31, 96, 31, 219, 31, 12, 31, 136, 31, 3, 31, 134, 31, 95, 31, 85, 31, 26, 31, 176, 31, 129, 31, 164, 31, 160, 31, 252, 31, 66, 31, 148, 31, 51, 31, 208, 31, 4, 31, 4, 30, 4, 29, 4, 28, 4, 27, 4, 26, 4, 25, 4, 24, 4, 23, 4, 22, 4, 21, 4, 20, 4, 19, 4, 18, 4, 17, 4, 16, 4, 15, 4, 14, 4, 13, 4, 12, 4, 11, 4, 10, 4, 9, 4, 8, 4, 7, 4, 6, 4, 5, 4, 4, 4, 3, 4, 2, 4, 1, 4, 0, 4, 0, 100, 31, 2, 31, 131, 31, 242, 31, 77, 31, 192, 31, 85, 31, 166, 31, 105, 31, 126, 31, 10, 31, 53, 31, 93, 31, 193, 31, 162, 31, 79, 31, 160, 31, 221, 31, 214, 31, 235, 31, 69, 31, 147, 31, 222, 31, 93, 31, 44, 31, 208, 31, 133, 31, 94, 31, 177, 31, 104, 31, 111, 31, 203, 31, 58, 31, 105, 31, 9, 31, 176, 31, 1, 31, 164, 31, 123, 31, 33, 31, 219, 31, 165, 31, 175, 31, 21, 31, 18, 31, 182, 31, 136, 31, 246, 31, 15, 31, 232, 31, 12, 31, 233, 31, 20, 31, 46, 31, 20, 31, 180, 31, 61, 31, 207, 31, 23, 31, 100, 31, 129, 31, 249, 31, 156, 31, 200, 31, 173, 31, 64, 31, 233, 31, 133, 31, 169, 31, 94, 31, 121, 31, 13, 31, 77, 31, 84, 31, 200, 31, 121, 31, 70, 31, 50, 31, 254, 31, 19, 31, 228, 31, 53, 31, 158, 31, 47, 31, 250, 31, 220, 31, 238, 31, 161, 31, 218, 31, 73, 31, 145, 31, 54, 31, 248, 31, 89, 31, 40, 31, 27, 31, 235, 31, 177, 31, 233, 31, 43, 31, 12, 31, 174, 31, 135, 31, 8, 31, 171, 31, 100, 31, 54, 31, 195, 31, 250, 31, 96, 31, 25, 31, 189, 31, 155, 31, 102, 31, 229, 31, 37, 31, 212, 31, 113, 31, 196, 31, 137, 31, 202, 31, 73, 31, 157, 31, 242, 31, 176, 31, 87, 31, 164, 31, 186, 31, 52, 31, 240, 31, 69, 31, 10, 31, 100, 31, 39, 31, 90, 31, 138, 31, 110, 31, 110, 30, 110, 29, 110, 28, 110, 27, 110, 26, 110, 25, 110, 24, 110, 23, 110, 22, 110, 21, 110, 20, 110, 19, 110, 18, 110, 17, 110, 16, 110, 15, 110, 14, 110, 13, 110, 12, 110, 11, 110, 10, 110, 9, 110, 8, 110, 7, 110, 6, 110, 5, 110, 4, 110, 3, 110, 2, 110, 1, 110, 0, 110, 0, 110, 0, 110, 0, 110, 0, 110, 0, 110, 0, 110, 0, 110, 0, 186, 31, 246, 31, 254, 31, 127, 31, 195, 31, 71, 31, 197, 31, 235, 31, 125, 31, 8, 31, 2, 31, 201, 31, 94, 31, 228, 31, 124, 31, 230, 31, 56, 31, 111, 31, 158, 31, 48, 31, 132, 31, 144, 31, 6, 31, 128, 31, 171, 31, 200, 31, 187, 31, 80, 31, 68, 31, 54, 31, 125, 31, 104, 31, 131, 31, 126, 31, 224, 31, 178, 31, 54, 31, 143, 31, 206, 31, 16, 31, 227, 31, 164, 31, 38, 31, 41, 31, 165, 31, 55, 31, 251, 31, 73, 31, 169, 31, 187, 31, 198, 31, 194, 31, 72, 31, 183, 31, 123, 31, 240, 31, 198, 31, 198, 30, 198, 29, 198, 28, 198, 27, 198, 26, 198, 25, 198, 24, 198, 23, 198, 22, 198, 21, 198, 20, 198, 19, 198, 18, 198, 17, 198, 16, 198, 15, 198, 14, 198, 13, 198, 12, 198, 11, 198, 10, 198, 9, 198, 8, 198, 7, 198, 6, 198, 5, 198, 4, 198, 3, 198, 2, 198, 1, 198, 0, 198, 0, 198, 0, 198, 0, 150, 31, 44, 31, 35, 31, 226, 31, 29, 31, 100, 31, 128, 31, 76, 31, 198, 31, 201, 31, 121, 31, 99, 31, 116, 31, 203, 31, 144, 31, 18, 31, 248, 31, 203, 31, 6, 31, 132, 31, 124, 31, 139, 31, 22, 31, 28, 31, 28, 30, 173, 31, 215, 31, 64, 31, 201, 31, 184, 31, 90, 31, 69, 31, 60, 31, 81, 31, 18, 31, 38, 31, 167, 31, 79, 31, 28, 31, 222, 31, 85, 31, 69, 31, 239, 31, 73, 31, 224, 31, 38, 31, 179, 31, 198, 31, 244, 31, 62, 31, 227, 31, 193, 31, 30, 31, 28, 31, 68, 31, 15, 31, 4, 31, 128, 31, 79, 31, 247, 31, 54, 31, 215, 31, 39, 31, 198, 31, 198, 30, 198, 29, 198, 28, 198, 27, 198, 26, 198, 25, 198, 24, 198, 23, 198, 22, 198, 21, 198, 20, 198, 19, 198, 18, 198, 17, 198, 16, 198, 15, 198, 14, 198, 13, 121, 31, 168, 31, 105, 31, 73, 31, 53, 31, 210, 31, 71, 31, 157, 31, 229, 31, 98, 31, 117, 31, 247, 31, 241, 31, 43, 31, 156, 31, 139, 31, 81, 31, 46, 31, 54, 31, 129, 31, 90, 31, 27, 31, 250, 31, 247, 31, 146, 31, 202, 31, 119, 31, 227, 31, 5, 31, 67, 31, 145, 31, 237, 31, 12, 31, 144, 31, 40, 31, 153, 31, 223, 31, 129, 31, 155, 31, 26, 31, 233, 31, 255, 31, 205, 31, 79, 31, 48, 31, 168, 31, 63, 31, 73, 31, 154, 31, 130, 31, 162, 31, 64, 31, 84, 31, 72, 31, 124, 31, 73, 31, 155, 31, 33, 31, 51, 31, 209, 31, 119, 31, 204, 31, 58, 31, 41, 31);
    constant SCENARIO_ADDRESS_2 : integer := 30012;


    -- third run

    constant SCENARIO_LENGTH_3 : integer := 628;
    type scenario_type_3 is array (0 to SCENARIO_LENGTH_3*2-1) of integer;
    signal scenario_input_3 : scenario_type_3 := (52, 0, 54, 0, 12, 0, 233, 0, 3, 0, 116, 0, 175, 0, 75, 0, 68, 0, 107, 0, 108, 0, 62, 0, 41, 0, 196, 0, 206, 0, 67, 0, 116, 0, 242, 0, 164, 0, 171, 0, 245, 0, 10, 0, 16, 0, 9, 0, 173, 0, 255, 0, 196, 0, 37, 0, 184, 0, 131, 0, 56, 0, 77, 0, 190, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 202, 0, 177, 0, 59, 0, 116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 0, 101, 0, 212, 0, 56, 0, 54, 0, 30, 0, 216, 0, 158, 0, 187, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 129, 0, 126, 0, 98, 0, 86, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 153, 0, 87, 0, 176, 0, 137, 0, 61, 0, 57, 0, 234, 0, 116, 0, 152, 0, 114, 0, 60, 0, 141, 0, 168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 190, 0, 60, 0, 141, 0, 53, 0, 53, 0, 206, 0, 176, 0, 200, 0, 77, 0, 16, 0, 194, 0, 89, 0, 171, 0, 105, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 206, 0, 124, 0, 117, 0, 187, 0, 62, 0, 218, 0, 236, 0, 145, 0, 71, 0, 50, 0, 248, 0, 236, 0, 18, 0, 219, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 208, 0, 94, 0, 221, 0, 205, 0, 239, 0, 241, 0, 116, 0, 63, 0, 122, 0, 75, 0, 29, 0, 249, 0, 12, 0, 17, 0, 71, 0, 190, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 189, 0, 203, 0, 41, 0, 76, 0, 21, 0, 170, 0, 100, 0, 230, 0, 37, 0, 177, 0, 214, 0, 208, 0, 250, 0, 112, 0, 100, 0, 201, 0, 137, 0, 219, 0, 125, 0, 98, 0, 12, 0, 123, 0, 39, 0, 63, 0, 117, 0, 176, 0, 100, 0, 106, 0, 24, 0, 227, 0, 206, 0, 55, 0, 82, 0, 1, 0, 153, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 0, 145, 0, 112, 0, 128, 0, 105, 0, 176, 0, 173, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 172, 0, 133, 0, 185, 0, 0, 0, 238, 0, 166, 0, 142, 0, 72, 0, 188, 0, 113, 0, 100, 0, 51, 0, 58, 0, 60, 0, 59, 0, 252, 0, 90, 0, 252, 0, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 0, 207, 0, 218, 0, 190, 0, 203, 0, 215, 0, 87, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);
    signal scenario_full_3  : scenario_type_3 := (52, 31, 54, 31, 12, 31, 233, 31, 3, 31, 116, 31, 175, 31, 75, 31, 68, 31, 107, 31, 108, 31, 62, 31, 41, 31, 196, 31, 206, 31, 67, 31, 116, 31, 242, 31, 164, 31, 171, 31, 245, 31, 10, 31, 16, 31, 9, 31, 173, 31, 255, 31, 196, 31, 37, 31, 184, 31, 131, 31, 56, 31, 77, 31, 190, 31, 60, 31, 60, 30, 60, 29, 60, 28, 60, 27, 60, 26, 60, 25, 60, 24, 60, 23, 60, 22, 60, 21, 60, 20, 60, 19, 60, 18, 60, 17, 60, 16, 60, 15, 60, 14, 60, 13, 60, 12, 60, 11, 60, 10, 60, 9, 60, 8, 60, 7, 60, 6, 60, 5, 60, 4, 60, 3, 60, 2, 60, 1, 202, 31, 177, 31, 59, 31, 116, 31, 116, 30, 116, 29, 116, 28, 116, 27, 116, 26, 116, 25, 116, 24, 116, 23, 116, 22, 116, 21, 116, 20, 116, 19, 116, 18, 116, 17, 116, 16, 116, 15, 116, 14, 116, 13, 116, 12, 116, 11, 116, 10, 116, 9, 116, 8, 116, 7, 116, 6, 116, 5, 116, 4, 116, 3, 116, 2, 116, 1, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 116, 0, 59, 31, 101, 31, 212, 31, 56, 31, 54, 31, 30, 31, 216, 31, 158, 31, 187, 31, 187, 30, 187, 29, 187, 28, 187, 27, 187, 26, 187, 25, 187, 24, 187, 23, 187, 22, 187, 21, 187, 20, 187, 19, 187, 18, 187, 17, 187, 16, 187, 15, 187, 14, 187, 13, 129, 31, 126, 31, 98, 31, 86, 31, 86, 30, 86, 29, 86, 28, 86, 27, 86, 26, 86, 25, 86, 24, 86, 23, 86, 22, 86, 21, 86, 20, 86, 19, 86, 18, 86, 17, 86, 16, 86, 15, 86, 14, 86, 13, 86, 12, 86, 11, 86, 10, 86, 9, 86, 8, 86, 7, 86, 6, 86, 5, 86, 4, 86, 3, 86, 2, 86, 1, 86, 0, 86, 0, 86, 0, 86, 0, 86, 0, 86, 0, 86, 0, 86, 0, 86, 0, 86, 0, 86, 0, 64, 31, 153, 31, 87, 31, 176, 31, 137, 31, 61, 31, 57, 31, 234, 31, 116, 31, 152, 31, 114, 31, 60, 31, 141, 31, 168, 31, 168, 30, 168, 29, 168, 28, 168, 27, 168, 26, 168, 25, 168, 24, 168, 23, 168, 22, 168, 21, 168, 20, 168, 19, 168, 18, 168, 17, 168, 16, 168, 15, 168, 14, 168, 13, 168, 12, 168, 11, 168, 10, 168, 9, 168, 8, 168, 7, 168, 6, 168, 5, 168, 4, 168, 3, 168, 2, 168, 1, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 168, 0, 190, 31, 60, 31, 141, 31, 53, 31, 53, 31, 206, 31, 176, 31, 200, 31, 77, 31, 16, 31, 194, 31, 89, 31, 171, 31, 105, 31, 105, 30, 105, 29, 105, 28, 105, 27, 105, 26, 105, 25, 105, 24, 105, 23, 105, 22, 105, 21, 105, 20, 105, 19, 105, 18, 105, 17, 105, 16, 105, 15, 105, 14, 105, 13, 105, 12, 105, 11, 105, 10, 105, 9, 105, 8, 105, 7, 105, 6, 105, 5, 105, 4, 105, 3, 105, 2, 105, 1, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 105, 0, 206, 31, 124, 31, 117, 31, 187, 31, 62, 31, 218, 31, 236, 31, 145, 31, 71, 31, 50, 31, 248, 31, 236, 31, 18, 31, 219, 31, 219, 30, 219, 29, 219, 28, 219, 27, 219, 26, 219, 25, 219, 24, 219, 23, 219, 22, 219, 21, 219, 20, 219, 19, 219, 18, 219, 17, 219, 16, 219, 15, 219, 14, 219, 13, 219, 12, 219, 11, 219, 10, 219, 9, 219, 8, 219, 7, 219, 6, 219, 5, 208, 31, 94, 31, 221, 31, 205, 31, 239, 31, 241, 31, 116, 31, 63, 31, 122, 31, 75, 31, 29, 31, 249, 31, 12, 31, 17, 31, 71, 31, 190, 31, 190, 30, 190, 29, 190, 28, 190, 27, 190, 26, 190, 25, 190, 24, 190, 23, 190, 22, 190, 21, 190, 20, 190, 19, 190, 18, 190, 17, 190, 16, 190, 15, 190, 14, 190, 13, 190, 12, 190, 11, 190, 10, 190, 9, 190, 8, 190, 7, 190, 6, 190, 5, 190, 4, 190, 3, 190, 2, 190, 1, 190, 0, 190, 0, 190, 0, 190, 0, 190, 0, 190, 0, 189, 31, 203, 31, 41, 31, 76, 31, 21, 31, 170, 31, 100, 31, 230, 31, 37, 31, 177, 31, 214, 31, 208, 31, 250, 31, 112, 31, 100, 31, 201, 31, 137, 31, 219, 31, 125, 31, 98, 31, 12, 31, 123, 31, 39, 31, 63, 31, 117, 31, 176, 31, 100, 31, 106, 31, 24, 31, 227, 31, 206, 31, 55, 31, 82, 31, 1, 31, 153, 31, 153, 30, 153, 29, 153, 28, 153, 27, 153, 26, 153, 25, 153, 24, 153, 23, 153, 22, 153, 21, 153, 20, 153, 19, 80, 31, 145, 31, 112, 31, 128, 31, 105, 31, 176, 31, 173, 31, 20, 31, 20, 30, 20, 29, 20, 28, 20, 27, 20, 26, 20, 25, 20, 24, 20, 23, 20, 22, 20, 21, 20, 20, 20, 19, 20, 18, 20, 17, 20, 16, 20, 15, 20, 14, 20, 13, 20, 12, 20, 11, 20, 10, 20, 9, 20, 8, 20, 7, 20, 6, 20, 5, 20, 4, 20, 3, 20, 2, 20, 1, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 20, 0, 13, 31, 172, 31, 133, 31, 185, 31, 185, 30, 238, 31, 166, 31, 142, 31, 72, 31, 188, 31, 113, 31, 100, 31, 51, 31, 58, 31, 60, 31, 59, 31, 252, 31, 90, 31, 252, 31, 68, 31, 68, 30, 68, 29, 68, 28, 68, 27, 68, 26, 68, 25, 68, 24, 68, 23, 68, 22, 68, 21, 68, 20, 68, 19, 68, 18, 68, 17, 68, 16, 68, 15, 68, 14, 68, 13, 68, 12, 68, 11, 68, 10, 68, 9, 68, 8, 68, 7, 68, 6, 68, 5, 68, 4, 68, 3, 68, 2, 80, 31, 207, 31, 218, 31, 190, 31, 203, 31, 215, 31, 87, 31, 33, 31, 33, 30, 33, 29, 33, 28, 33, 27, 33, 26, 33, 25, 33, 24, 33, 23, 33, 22, 33, 21, 33, 20, 33, 19, 33, 18, 33, 17, 33, 16, 33, 15, 33, 14, 33, 13, 33, 12, 33, 11, 33, 10, 33, 9, 33, 8, 33, 7, 33, 6, 33, 5, 33, 4, 33, 3, 33, 2, 33, 1, 33, 31, 78, 31, 78, 30, 78, 29, 78, 28, 78, 27, 78, 26, 78, 25, 78, 24, 78, 23);
    constant SCENARIO_ADDRESS_3 : integer := 40000;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;


        -- Configure second run
        
        for i in 0 to SCENARIO_LENGTH_2*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_2+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_2(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        -- Configure third run

        for i in 0 to SCENARIO_LENGTH_3*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_3+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input_3(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';

        -- start sencond run without reset

        wait for 50 ns;

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_2, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_2, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';

        -- start third run without reset

        wait for 50 ns;

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS_3, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH_3, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
        
        wait for 5 ns;
        
        tb_start <= '0';

        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);


        -- second run
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH_2*2-1 loop
            assert RAM(SCENARIO_ADDRESS_2+i) = std_logic_vector(to_unsigned(scenario_full_2(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_2(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);



        -- third run
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH_3*2-1 loop
            assert RAM(SCENARIO_ADDRESS_3+i) = std_logic_vector(to_unsigned(scenario_full_3(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full_3(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);



        -- end

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
